// +FHDR -----------------------------------------------------------------------
// Copyright (c) Silicon Optronics. Inc. 2022
//
// File Name:           cube root lut 
// Author:              Willy Lin
// Version:             1.0
// Date:                2022/10/25
// Last Modified On:
// Last Modified By:    $Author$
//
// File precision  : input  : 8.4
//                   output : 0~1     : 0.14
//                            1~8     : 1.13
//                            8~64    : 2.12
//                            64~256  : 3.11
//
// -FHDR -----------------------------------------------------------------------

module cube_lut_12_14_ver2
(
//----------------------------------------------//
// Output declaration                           //
//----------------------------------------------//
    output reg [13:0] o_data,
    output reg [1:0]  o_prcis_idx,
//----------------------------------------------//
// Input declaration                            //
//----------------------------------------------//
    input      [11:0] i_data,
    input             clk,
    input             rst_n
);

//----------------------------------------------//
// Local Parameter                              //
//----------------------------------------------//

//----------------------------------------------//
// Register & Wire declaration                  //
//----------------------------------------------//
wire        decode_0;
wire        decode_1;
wire        decode_2;
wire        decode_3;
wire        decode_4;
wire        decode_5;
wire        decode_6;
wire        decode_7;

wire [13:0] com_lut;

reg  [13:0] cube_lut_0;
reg  [13:0] cube_lut_1;
reg  [13:0] cube_lut_2;
reg  [13:0] cube_lut_3;
reg  [13:0] cube_lut_4;
reg  [13:0] cube_lut_5;
reg  [13:0] cube_lut_6;
reg  [13:0] cube_lut_7;

//output port 
wire [1:0]  o_prcis_idx_nxt;
wire [13:0] o_data_nxt;

//----------------------------------------------//
// Code Descriptions                            //
//----------------------------------------------//
//find region 
assign o_prcis_idx_nxt  = (i_data[11:4] <8) ? (i_data[11:4] <1)  ? 2'b00 : 2'b01 : 
                                              (i_data[11:4] <64) ? 2'b10 : 2'b11 ;


assign decode_0         = i_data[11:9] == 3'b000;
assign decode_1         = i_data[11:9] == 3'b001;
assign decode_2         = i_data[11:9] == 3'b010;
assign decode_3         = i_data[11:9] == 3'b011;
assign decode_4         = i_data[11:9] == 3'b100;
assign decode_5         = i_data[11:9] == 3'b101;
assign decode_6         = i_data[11:9] == 3'b110;
assign decode_7         = i_data[11:9] == 3'b111;

assign com_lut          = ({14{decode_0}} & cube_lut_0) |
                          ({14{decode_1}} & cube_lut_1) |
                          ({14{decode_2}} & cube_lut_2) |
                          ({14{decode_3}} & cube_lut_3) |
                          ({14{decode_4}} & cube_lut_4) |
                          ({14{decode_5}} & cube_lut_5) |
                          ({14{decode_6}} & cube_lut_6) |
                          ({14{decode_7}} & cube_lut_7);

assign o_data_nxt       = com_lut;

always@* begin
    
    cube_lut_0 = 0;
    
    case(i_data[8:0])
 
 9'd0   : cube_lut_0 = 14'b0;
9'd1   : cube_lut_0 = 14'b01100101100101;
9'd2   : cube_lut_0 = 14'b10000000000000;
9'd3   : cube_lut_0 = 14'b10010010100001;
9'd4   : cube_lut_0 = 14'b10100001010001;
9'd5   : cube_lut_0 = 14'b10101101101110;
9'd6   : cube_lut_0 = 14'b10111000100110;
9'd7   : cube_lut_0 = 14'b11000010010101;
9'd8   : cube_lut_0 = 14'b11001011001011;
9'd9   : cube_lut_0 = 14'b11010011010100;
9'd10   : cube_lut_0 = 14'b11011010111000;
9'd11   : cube_lut_0 = 14'b11100001111100;
9'd12   : cube_lut_0 = 14'b11101000100101;
9'd13   : cube_lut_0 = 14'b11101110111000;
9'd14   : cube_lut_0 = 14'b11110100110110;
9'd15   : cube_lut_0 = 14'b11111010100011;
9'd16   : cube_lut_0 = 14'b10000000000000;
9'd17   : cube_lut_0 = 14'b10000010100111;
9'd18   : cube_lut_0 = 14'b10000101001000;
9'd19   : cube_lut_0 = 14'b10000111100010;
9'd20   : cube_lut_0 = 14'b10001001111000;
9'd21   : cube_lut_0 = 14'b10001100001001;
9'd22   : cube_lut_0 = 14'b10001110010101;
9'd23   : cube_lut_0 = 14'b10010000011101;
9'd24   : cube_lut_0 = 14'b10010010100001;
9'd25   : cube_lut_0 = 14'b10010100100001;
9'd26   : cube_lut_0 = 14'b10010110011111;
9'd27   : cube_lut_0 = 14'b10011000011000;
9'd28   : cube_lut_0 = 14'b10011010001111;
9'd29   : cube_lut_0 = 14'b10011100000100;
9'd30   : cube_lut_0 = 14'b10011101110101;
9'd31   : cube_lut_0 = 14'b10011111100100;
9'd32   : cube_lut_0 = 14'b10100001010001;
9'd33   : cube_lut_0 = 14'b10100010111011;
9'd34   : cube_lut_0 = 14'b10100100100011;
9'd35   : cube_lut_0 = 14'b10100110001010;
9'd36   : cube_lut_0 = 14'b10100111101110;
9'd37   : cube_lut_0 = 14'b10101001010001;
9'd38   : cube_lut_0 = 14'b10101010110001;
9'd39   : cube_lut_0 = 14'b10101100010000;
9'd40   : cube_lut_0 = 14'b10101101101110;
9'd41   : cube_lut_0 = 14'b10101111001010;
9'd42   : cube_lut_0 = 14'b10110000100100;
9'd43   : cube_lut_0 = 14'b10110001111101;
9'd44   : cube_lut_0 = 14'b10110011010101;
9'd45   : cube_lut_0 = 14'b10110100101011;
9'd46   : cube_lut_0 = 14'b10110110000000;
9'd47   : cube_lut_0 = 14'b10110111010100;
9'd48   : cube_lut_0 = 14'b10111000100110;
9'd49   : cube_lut_0 = 14'b10111001111000;
9'd50   : cube_lut_0 = 14'b10111011001000;
9'd51   : cube_lut_0 = 14'b10111100011000;
9'd52   : cube_lut_0 = 14'b10111101100110;
9'd53   : cube_lut_0 = 14'b10111110110011;
9'd54   : cube_lut_0 = 14'b11000000000000;
9'd55   : cube_lut_0 = 14'b11000001001011;
9'd56   : cube_lut_0 = 14'b11000010010101;
9'd57   : cube_lut_0 = 14'b11000011011111;
9'd58   : cube_lut_0 = 14'b11000100101000;
9'd59   : cube_lut_0 = 14'b11000101110000;
9'd60   : cube_lut_0 = 14'b11000110110111;
9'd61   : cube_lut_0 = 14'b11000111111101;
9'd62   : cube_lut_0 = 14'b11001001000011;
9'd63   : cube_lut_0 = 14'b11001010000111;
9'd64   : cube_lut_0 = 14'b11001011001011;
9'd65   : cube_lut_0 = 14'b11001100001111;
9'd66   : cube_lut_0 = 14'b11001101010010;
9'd67   : cube_lut_0 = 14'b11001110010100;
9'd68   : cube_lut_0 = 14'b11001111010101;
9'd69   : cube_lut_0 = 14'b11010000010110;
9'd70   : cube_lut_0 = 14'b11010001010110;
9'd71   : cube_lut_0 = 14'b11010010010101;
9'd72   : cube_lut_0 = 14'b11010011010100;
9'd73   : cube_lut_0 = 14'b11010100010011;
9'd74   : cube_lut_0 = 14'b11010101010000;
9'd75   : cube_lut_0 = 14'b11010110001101;
9'd76   : cube_lut_0 = 14'b11010111001010;
9'd77   : cube_lut_0 = 14'b11011000000110;
9'd78   : cube_lut_0 = 14'b11011001000010;
9'd79   : cube_lut_0 = 14'b11011001111101;
9'd80   : cube_lut_0 = 14'b11011010111000;
9'd81   : cube_lut_0 = 14'b11011011110010;
9'd82   : cube_lut_0 = 14'b11011100101011;
9'd83   : cube_lut_0 = 14'b11011101100101;
9'd84   : cube_lut_0 = 14'b11011110011101;
9'd85   : cube_lut_0 = 14'b11011111010110;
9'd86   : cube_lut_0 = 14'b11100000001101;
9'd87   : cube_lut_0 = 14'b11100001000101;
9'd88   : cube_lut_0 = 14'b11100001111100;
9'd89   : cube_lut_0 = 14'b11100010110010;
9'd90   : cube_lut_0 = 14'b11100011101001;
9'd91   : cube_lut_0 = 14'b11100100011110;
9'd92   : cube_lut_0 = 14'b11100101010100;
9'd93   : cube_lut_0 = 14'b11100110001001;
9'd94   : cube_lut_0 = 14'b11100110111101;
9'd95   : cube_lut_0 = 14'b11100111110001;
9'd96   : cube_lut_0 = 14'b11101000100101;
9'd97   : cube_lut_0 = 14'b11101001011001;
9'd98   : cube_lut_0 = 14'b11101010001100;
9'd99   : cube_lut_0 = 14'b11101010111111;
9'd100   : cube_lut_0 = 14'b11101011110001;
9'd101   : cube_lut_0 = 14'b11101100100011;
9'd102   : cube_lut_0 = 14'b11101101010101;
9'd103   : cube_lut_0 = 14'b11101110000111;
9'd104   : cube_lut_0 = 14'b11101110111000;
9'd105   : cube_lut_0 = 14'b11101111101001;
9'd106   : cube_lut_0 = 14'b11110000011001;
9'd107   : cube_lut_0 = 14'b11110001001001;
9'd108   : cube_lut_0 = 14'b11110001111001;
9'd109   : cube_lut_0 = 14'b11110010101001;
9'd110   : cube_lut_0 = 14'b11110011011000;
9'd111   : cube_lut_0 = 14'b11110100000111;
9'd112   : cube_lut_0 = 14'b11110100110110;
9'd113   : cube_lut_0 = 14'b11110101100101;
9'd114   : cube_lut_0 = 14'b11110110010011;
9'd115   : cube_lut_0 = 14'b11110111000001;
9'd116   : cube_lut_0 = 14'b11110111101111;
9'd117   : cube_lut_0 = 14'b11111000011100;
9'd118   : cube_lut_0 = 14'b11111001001001;
9'd119   : cube_lut_0 = 14'b11111001110110;
9'd120   : cube_lut_0 = 14'b11111010100011;
9'd121   : cube_lut_0 = 14'b11111011001111;
9'd122   : cube_lut_0 = 14'b11111011111011;
9'd123   : cube_lut_0 = 14'b11111100100111;
9'd124   : cube_lut_0 = 14'b11111101010011;
9'd125   : cube_lut_0 = 14'b11111101111110;
9'd126   : cube_lut_0 = 14'b11111110101010;
9'd127   : cube_lut_0 = 14'b11111111010101;
9'd128   : cube_lut_0 = 14'b10000000000000;
9'd129   : cube_lut_0 = 14'b10000000010101;
9'd130   : cube_lut_0 = 14'b10000000101010;
9'd131   : cube_lut_0 = 14'b10000000111111;
9'd132   : cube_lut_0 = 14'b10000001010100;
9'd133   : cube_lut_0 = 14'b10000001101001;
9'd134   : cube_lut_0 = 14'b10000001111110;
9'd135   : cube_lut_0 = 14'b10000010010010;
9'd136   : cube_lut_0 = 14'b10000010100111;
9'd137   : cube_lut_0 = 14'b10000010111011;
9'd138   : cube_lut_0 = 14'b10000011010000;
9'd139   : cube_lut_0 = 14'b10000011100100;
9'd140   : cube_lut_0 = 14'b10000011111000;
9'd141   : cube_lut_0 = 14'b10000100001100;
9'd142   : cube_lut_0 = 14'b10000100100000;
9'd143   : cube_lut_0 = 14'b10000100110100;
9'd144   : cube_lut_0 = 14'b10000101001000;
9'd145   : cube_lut_0 = 14'b10000101011011;
9'd146   : cube_lut_0 = 14'b10000101101111;
9'd147   : cube_lut_0 = 14'b10000110000010;
9'd148   : cube_lut_0 = 14'b10000110010110;
9'd149   : cube_lut_0 = 14'b10000110101001;
9'd150   : cube_lut_0 = 14'b10000110111100;
9'd151   : cube_lut_0 = 14'b10000111001111;
9'd152   : cube_lut_0 = 14'b10000111100010;
9'd153   : cube_lut_0 = 14'b10000111110101;
9'd154   : cube_lut_0 = 14'b10001000001000;
9'd155   : cube_lut_0 = 14'b10001000011011;
9'd156   : cube_lut_0 = 14'b10001000101110;
9'd157   : cube_lut_0 = 14'b10001001000001;
9'd158   : cube_lut_0 = 14'b10001001010011;
9'd159   : cube_lut_0 = 14'b10001001100110;
9'd160   : cube_lut_0 = 14'b10001001111000;
9'd161   : cube_lut_0 = 14'b10001010001010;
9'd162   : cube_lut_0 = 14'b10001010011101;
9'd163   : cube_lut_0 = 14'b10001010101111;
9'd164   : cube_lut_0 = 14'b10001011000001;
9'd165   : cube_lut_0 = 14'b10001011010011;
9'd166   : cube_lut_0 = 14'b10001011100101;
9'd167   : cube_lut_0 = 14'b10001011110111;
9'd168   : cube_lut_0 = 14'b10001100001001;
9'd169   : cube_lut_0 = 14'b10001100011011;
9'd170   : cube_lut_0 = 14'b10001100101100;
9'd171   : cube_lut_0 = 14'b10001100111110;
9'd172   : cube_lut_0 = 14'b10001101001111;
9'd173   : cube_lut_0 = 14'b10001101100001;
9'd174   : cube_lut_0 = 14'b10001101110010;
9'd175   : cube_lut_0 = 14'b10001110000100;
9'd176   : cube_lut_0 = 14'b10001110010101;
9'd177   : cube_lut_0 = 14'b10001110100110;
9'd178   : cube_lut_0 = 14'b10001110110111;
9'd179   : cube_lut_0 = 14'b10001111001000;
9'd180   : cube_lut_0 = 14'b10001111011001;
9'd181   : cube_lut_0 = 14'b10001111101010;
9'd182   : cube_lut_0 = 14'b10001111111011;
9'd183   : cube_lut_0 = 14'b10010000001100;
9'd184   : cube_lut_0 = 14'b10010000011101;
9'd185   : cube_lut_0 = 14'b10010000101110;
9'd186   : cube_lut_0 = 14'b10010000111110;
9'd187   : cube_lut_0 = 14'b10010001001111;
9'd188   : cube_lut_0 = 14'b10010001011111;
9'd189   : cube_lut_0 = 14'b10010001110000;
9'd190   : cube_lut_0 = 14'b10010010000000;
9'd191   : cube_lut_0 = 14'b10010010010001;
9'd192   : cube_lut_0 = 14'b10010010100001;
9'd193   : cube_lut_0 = 14'b10010010110001;
9'd194   : cube_lut_0 = 14'b10010011000001;
9'd195   : cube_lut_0 = 14'b10010011010010;
9'd196   : cube_lut_0 = 14'b10010011100010;
9'd197   : cube_lut_0 = 14'b10010011110010;
9'd198   : cube_lut_0 = 14'b10010100000010;
9'd199   : cube_lut_0 = 14'b10010100010010;
9'd200   : cube_lut_0 = 14'b10010100100001;
9'd201   : cube_lut_0 = 14'b10010100110001;
9'd202   : cube_lut_0 = 14'b10010101000001;
9'd203   : cube_lut_0 = 14'b10010101010001;
9'd204   : cube_lut_0 = 14'b10010101100000;
9'd205   : cube_lut_0 = 14'b10010101110000;
9'd206   : cube_lut_0 = 14'b10010110000000;
9'd207   : cube_lut_0 = 14'b10010110001111;
9'd208   : cube_lut_0 = 14'b10010110011111;
9'd209   : cube_lut_0 = 14'b10010110101110;
9'd210   : cube_lut_0 = 14'b10010110111101;
9'd211   : cube_lut_0 = 14'b10010111001101;
9'd212   : cube_lut_0 = 14'b10010111011100;
9'd213   : cube_lut_0 = 14'b10010111101011;
9'd214   : cube_lut_0 = 14'b10010111111010;
9'd215   : cube_lut_0 = 14'b10011000001001;
9'd216   : cube_lut_0 = 14'b10011000011000;
9'd217   : cube_lut_0 = 14'b10011000101000;
9'd218   : cube_lut_0 = 14'b10011000110111;
9'd219   : cube_lut_0 = 14'b10011001000101;
9'd220   : cube_lut_0 = 14'b10011001010100;
9'd221   : cube_lut_0 = 14'b10011001100011;
9'd222   : cube_lut_0 = 14'b10011001110010;
9'd223   : cube_lut_0 = 14'b10011010000001;
9'd224   : cube_lut_0 = 14'b10011010001111;
9'd225   : cube_lut_0 = 14'b10011010011110;
9'd226   : cube_lut_0 = 14'b10011010101101;
9'd227   : cube_lut_0 = 14'b10011010111011;
9'd228   : cube_lut_0 = 14'b10011011001010;
9'd229   : cube_lut_0 = 14'b10011011011000;
9'd230   : cube_lut_0 = 14'b10011011100111;
9'd231   : cube_lut_0 = 14'b10011011110101;
9'd232   : cube_lut_0 = 14'b10011100000100;
9'd233   : cube_lut_0 = 14'b10011100010010;
9'd234   : cube_lut_0 = 14'b10011100100000;
9'd235   : cube_lut_0 = 14'b10011100101110;
9'd236   : cube_lut_0 = 14'b10011100111101;
9'd237   : cube_lut_0 = 14'b10011101001011;
9'd238   : cube_lut_0 = 14'b10011101011001;
9'd239   : cube_lut_0 = 14'b10011101100111;
9'd240   : cube_lut_0 = 14'b10011101110101;
9'd241   : cube_lut_0 = 14'b10011110000011;
9'd242   : cube_lut_0 = 14'b10011110010001;
9'd243   : cube_lut_0 = 14'b10011110011111;
9'd244   : cube_lut_0 = 14'b10011110101101;
9'd245   : cube_lut_0 = 14'b10011110111011;
9'd246   : cube_lut_0 = 14'b10011111001001;
9'd247   : cube_lut_0 = 14'b10011111010110;
9'd248   : cube_lut_0 = 14'b10011111100100;
9'd249   : cube_lut_0 = 14'b10011111110010;
9'd250   : cube_lut_0 = 14'b10100000000000;
9'd251   : cube_lut_0 = 14'b10100000001101;
9'd252   : cube_lut_0 = 14'b10100000011011;
9'd253   : cube_lut_0 = 14'b10100000101000;
9'd254   : cube_lut_0 = 14'b10100000110110;
9'd255   : cube_lut_0 = 14'b10100001000011;
9'd256   : cube_lut_0 = 14'b10100001010001;
9'd257   : cube_lut_0 = 14'b10100001011110;
9'd258   : cube_lut_0 = 14'b10100001101100;
9'd259   : cube_lut_0 = 14'b10100001111001;
9'd260   : cube_lut_0 = 14'b10100010000110;
9'd261   : cube_lut_0 = 14'b10100010010100;
9'd262   : cube_lut_0 = 14'b10100010100001;
9'd263   : cube_lut_0 = 14'b10100010101110;
9'd264   : cube_lut_0 = 14'b10100010111011;
9'd265   : cube_lut_0 = 14'b10100011001000;
9'd266   : cube_lut_0 = 14'b10100011010101;
9'd267   : cube_lut_0 = 14'b10100011100011;
9'd268   : cube_lut_0 = 14'b10100011110000;
9'd269   : cube_lut_0 = 14'b10100011111101;
9'd270   : cube_lut_0 = 14'b10100100001010;
9'd271   : cube_lut_0 = 14'b10100100010111;
9'd272   : cube_lut_0 = 14'b10100100100011;
9'd273   : cube_lut_0 = 14'b10100100110000;
9'd274   : cube_lut_0 = 14'b10100100111101;
9'd275   : cube_lut_0 = 14'b10100101001010;
9'd276   : cube_lut_0 = 14'b10100101010111;
9'd277   : cube_lut_0 = 14'b10100101100100;
9'd278   : cube_lut_0 = 14'b10100101110000;
9'd279   : cube_lut_0 = 14'b10100101111101;
9'd280   : cube_lut_0 = 14'b10100110001010;
9'd281   : cube_lut_0 = 14'b10100110010110;
9'd282   : cube_lut_0 = 14'b10100110100011;
9'd283   : cube_lut_0 = 14'b10100110110000;
9'd284   : cube_lut_0 = 14'b10100110111100;
9'd285   : cube_lut_0 = 14'b10100111001001;
9'd286   : cube_lut_0 = 14'b10100111010101;
9'd287   : cube_lut_0 = 14'b10100111100010;
9'd288   : cube_lut_0 = 14'b10100111101110;
9'd289   : cube_lut_0 = 14'b10100111111010;
9'd290   : cube_lut_0 = 14'b10101000000111;
9'd291   : cube_lut_0 = 14'b10101000010011;
9'd292   : cube_lut_0 = 14'b10101000100000;
9'd293   : cube_lut_0 = 14'b10101000101100;
9'd294   : cube_lut_0 = 14'b10101000111000;
9'd295   : cube_lut_0 = 14'b10101001000100;
9'd296   : cube_lut_0 = 14'b10101001010001;
9'd297   : cube_lut_0 = 14'b10101001011101;
9'd298   : cube_lut_0 = 14'b10101001101001;
9'd299   : cube_lut_0 = 14'b10101001110101;
9'd300   : cube_lut_0 = 14'b10101010000001;
9'd301   : cube_lut_0 = 14'b10101010001101;
9'd302   : cube_lut_0 = 14'b10101010011001;
9'd303   : cube_lut_0 = 14'b10101010100101;
9'd304   : cube_lut_0 = 14'b10101010110001;
9'd305   : cube_lut_0 = 14'b10101010111101;
9'd306   : cube_lut_0 = 14'b10101011001001;
9'd307   : cube_lut_0 = 14'b10101011010101;
9'd308   : cube_lut_0 = 14'b10101011100001;
9'd309   : cube_lut_0 = 14'b10101011101101;
9'd310   : cube_lut_0 = 14'b10101011111001;
9'd311   : cube_lut_0 = 14'b10101100000101;
9'd312   : cube_lut_0 = 14'b10101100010000;
9'd313   : cube_lut_0 = 14'b10101100011100;
9'd314   : cube_lut_0 = 14'b10101100101000;
9'd315   : cube_lut_0 = 14'b10101100110100;
9'd316   : cube_lut_0 = 14'b10101100111111;
9'd317   : cube_lut_0 = 14'b10101101001011;
9'd318   : cube_lut_0 = 14'b10101101010111;
9'd319   : cube_lut_0 = 14'b10101101100010;
9'd320   : cube_lut_0 = 14'b10101101101110;
9'd321   : cube_lut_0 = 14'b10101101111001;
9'd322   : cube_lut_0 = 14'b10101110000101;
9'd323   : cube_lut_0 = 14'b10101110010000;
9'd324   : cube_lut_0 = 14'b10101110011100;
9'd325   : cube_lut_0 = 14'b10101110100111;
9'd326   : cube_lut_0 = 14'b10101110110011;
9'd327   : cube_lut_0 = 14'b10101110111110;
9'd328   : cube_lut_0 = 14'b10101111001010;
9'd329   : cube_lut_0 = 14'b10101111010101;
9'd330   : cube_lut_0 = 14'b10101111100000;
9'd331   : cube_lut_0 = 14'b10101111101100;
9'd332   : cube_lut_0 = 14'b10101111110111;
9'd333   : cube_lut_0 = 14'b10110000000010;
9'd334   : cube_lut_0 = 14'b10110000001110;
9'd335   : cube_lut_0 = 14'b10110000011001;
9'd336   : cube_lut_0 = 14'b10110000100100;
9'd337   : cube_lut_0 = 14'b10110000101111;
9'd338   : cube_lut_0 = 14'b10110000111010;
9'd339   : cube_lut_0 = 14'b10110001000110;
9'd340   : cube_lut_0 = 14'b10110001010001;
9'd341   : cube_lut_0 = 14'b10110001011100;
9'd342   : cube_lut_0 = 14'b10110001100111;
9'd343   : cube_lut_0 = 14'b10110001110010;
9'd344   : cube_lut_0 = 14'b10110001111101;
9'd345   : cube_lut_0 = 14'b10110010001000;
9'd346   : cube_lut_0 = 14'b10110010010011;
9'd347   : cube_lut_0 = 14'b10110010011110;
9'd348   : cube_lut_0 = 14'b10110010101001;
9'd349   : cube_lut_0 = 14'b10110010110100;
9'd350   : cube_lut_0 = 14'b10110010111111;
9'd351   : cube_lut_0 = 14'b10110011001010;
9'd352   : cube_lut_0 = 14'b10110011010101;
9'd353   : cube_lut_0 = 14'b10110011100000;
9'd354   : cube_lut_0 = 14'b10110011101010;
9'd355   : cube_lut_0 = 14'b10110011110101;
9'd356   : cube_lut_0 = 14'b10110100000000;
9'd357   : cube_lut_0 = 14'b10110100001011;
9'd358   : cube_lut_0 = 14'b10110100010101;
9'd359   : cube_lut_0 = 14'b10110100100000;
9'd360   : cube_lut_0 = 14'b10110100101011;
9'd361   : cube_lut_0 = 14'b10110100110110;
9'd362   : cube_lut_0 = 14'b10110101000000;
9'd363   : cube_lut_0 = 14'b10110101001011;
9'd364   : cube_lut_0 = 14'b10110101010110;
9'd365   : cube_lut_0 = 14'b10110101100000;
9'd366   : cube_lut_0 = 14'b10110101101011;
9'd367   : cube_lut_0 = 14'b10110101110101;
9'd368   : cube_lut_0 = 14'b10110110000000;
9'd369   : cube_lut_0 = 14'b10110110001011;
9'd370   : cube_lut_0 = 14'b10110110010101;
9'd371   : cube_lut_0 = 14'b10110110100000;
9'd372   : cube_lut_0 = 14'b10110110101010;
9'd373   : cube_lut_0 = 14'b10110110110100;
9'd374   : cube_lut_0 = 14'b10110110111111;
9'd375   : cube_lut_0 = 14'b10110111001001;
9'd376   : cube_lut_0 = 14'b10110111010100;
9'd377   : cube_lut_0 = 14'b10110111011110;
9'd378   : cube_lut_0 = 14'b10110111101001;
9'd379   : cube_lut_0 = 14'b10110111110011;
9'd380   : cube_lut_0 = 14'b10110111111101;
9'd381   : cube_lut_0 = 14'b10111000001000;
9'd382   : cube_lut_0 = 14'b10111000010010;
9'd383   : cube_lut_0 = 14'b10111000011100;
9'd384   : cube_lut_0 = 14'b10111000100110;
9'd385   : cube_lut_0 = 14'b10111000110001;
9'd386   : cube_lut_0 = 14'b10111000111011;
9'd387   : cube_lut_0 = 14'b10111001000101;
9'd388   : cube_lut_0 = 14'b10111001001111;
9'd389   : cube_lut_0 = 14'b10111001011001;
9'd390   : cube_lut_0 = 14'b10111001100100;
9'd391   : cube_lut_0 = 14'b10111001101110;
9'd392   : cube_lut_0 = 14'b10111001111000;
9'd393   : cube_lut_0 = 14'b10111010000010;
9'd394   : cube_lut_0 = 14'b10111010001100;
9'd395   : cube_lut_0 = 14'b10111010010110;
9'd396   : cube_lut_0 = 14'b10111010100000;
9'd397   : cube_lut_0 = 14'b10111010101010;
9'd398   : cube_lut_0 = 14'b10111010110100;
9'd399   : cube_lut_0 = 14'b10111010111110;
9'd400   : cube_lut_0 = 14'b10111011001000;
9'd401   : cube_lut_0 = 14'b10111011010010;
9'd402   : cube_lut_0 = 14'b10111011011100;
9'd403   : cube_lut_0 = 14'b10111011100110;
9'd404   : cube_lut_0 = 14'b10111011110000;
9'd405   : cube_lut_0 = 14'b10111011111010;
9'd406   : cube_lut_0 = 14'b10111100000100;
9'd407   : cube_lut_0 = 14'b10111100001110;
9'd408   : cube_lut_0 = 14'b10111100011000;
9'd409   : cube_lut_0 = 14'b10111100100001;
9'd410   : cube_lut_0 = 14'b10111100101011;
9'd411   : cube_lut_0 = 14'b10111100110101;
9'd412   : cube_lut_0 = 14'b10111100111111;
9'd413   : cube_lut_0 = 14'b10111101001001;
9'd414   : cube_lut_0 = 14'b10111101010010;
9'd415   : cube_lut_0 = 14'b10111101011100;
9'd416   : cube_lut_0 = 14'b10111101100110;
9'd417   : cube_lut_0 = 14'b10111101110000;
9'd418   : cube_lut_0 = 14'b10111101111001;
9'd419   : cube_lut_0 = 14'b10111110000011;
9'd420   : cube_lut_0 = 14'b10111110001101;
9'd421   : cube_lut_0 = 14'b10111110010110;
9'd422   : cube_lut_0 = 14'b10111110100000;
9'd423   : cube_lut_0 = 14'b10111110101010;
9'd424   : cube_lut_0 = 14'b10111110110011;
9'd425   : cube_lut_0 = 14'b10111110111101;
9'd426   : cube_lut_0 = 14'b10111111000110;
9'd427   : cube_lut_0 = 14'b10111111010000;
9'd428   : cube_lut_0 = 14'b10111111011001;
9'd429   : cube_lut_0 = 14'b10111111100011;
9'd430   : cube_lut_0 = 14'b10111111101101;
9'd431   : cube_lut_0 = 14'b10111111110110;
9'd432   : cube_lut_0 = 14'b11000000000000;
9'd433   : cube_lut_0 = 14'b11000000001001;
9'd434   : cube_lut_0 = 14'b11000000010010;
9'd435   : cube_lut_0 = 14'b11000000011100;
9'd436   : cube_lut_0 = 14'b11000000100101;
9'd437   : cube_lut_0 = 14'b11000000101111;
9'd438   : cube_lut_0 = 14'b11000000111000;
9'd439   : cube_lut_0 = 14'b11000001000010;
9'd440   : cube_lut_0 = 14'b11000001001011;
9'd441   : cube_lut_0 = 14'b11000001010100;
9'd442   : cube_lut_0 = 14'b11000001011110;
9'd443   : cube_lut_0 = 14'b11000001100111;
9'd444   : cube_lut_0 = 14'b11000001110000;
9'd445   : cube_lut_0 = 14'b11000001111010;
9'd446   : cube_lut_0 = 14'b11000010000011;
9'd447   : cube_lut_0 = 14'b11000010001100;
9'd448   : cube_lut_0 = 14'b11000010010101;
9'd449   : cube_lut_0 = 14'b11000010011111;
9'd450   : cube_lut_0 = 14'b11000010101000;
9'd451   : cube_lut_0 = 14'b11000010110001;
9'd452   : cube_lut_0 = 14'b11000010111010;
9'd453   : cube_lut_0 = 14'b11000011000011;
9'd454   : cube_lut_0 = 14'b11000011001101;
9'd455   : cube_lut_0 = 14'b11000011010110;
9'd456   : cube_lut_0 = 14'b11000011011111;
9'd457   : cube_lut_0 = 14'b11000011101000;
9'd458   : cube_lut_0 = 14'b11000011110001;
9'd459   : cube_lut_0 = 14'b11000011111010;
9'd460   : cube_lut_0 = 14'b11000100000011;
9'd461   : cube_lut_0 = 14'b11000100001101;
9'd462   : cube_lut_0 = 14'b11000100010110;
9'd463   : cube_lut_0 = 14'b11000100011111;
9'd464   : cube_lut_0 = 14'b11000100101000;
9'd465   : cube_lut_0 = 14'b11000100110001;
9'd466   : cube_lut_0 = 14'b11000100111010;
9'd467   : cube_lut_0 = 14'b11000101000011;
9'd468   : cube_lut_0 = 14'b11000101001100;
9'd469   : cube_lut_0 = 14'b11000101010101;
9'd470   : cube_lut_0 = 14'b11000101011110;
9'd471   : cube_lut_0 = 14'b11000101100111;
9'd472   : cube_lut_0 = 14'b11000101110000;
9'd473   : cube_lut_0 = 14'b11000101111001;
9'd474   : cube_lut_0 = 14'b11000110000001;
9'd475   : cube_lut_0 = 14'b11000110001010;
9'd476   : cube_lut_0 = 14'b11000110010011;
9'd477   : cube_lut_0 = 14'b11000110011100;
9'd478   : cube_lut_0 = 14'b11000110100101;
9'd479   : cube_lut_0 = 14'b11000110101110;
9'd480   : cube_lut_0 = 14'b11000110110111;
9'd481   : cube_lut_0 = 14'b11000111000000;
9'd482   : cube_lut_0 = 14'b11000111001000;
9'd483   : cube_lut_0 = 14'b11000111010001;
9'd484   : cube_lut_0 = 14'b11000111011010;
9'd485   : cube_lut_0 = 14'b11000111100011;
9'd486   : cube_lut_0 = 14'b11000111101100;
9'd487   : cube_lut_0 = 14'b11000111110100;
9'd488   : cube_lut_0 = 14'b11000111111101;
9'd489   : cube_lut_0 = 14'b11001000000110;
9'd490   : cube_lut_0 = 14'b11001000001111;
9'd491   : cube_lut_0 = 14'b11001000010111;
9'd492   : cube_lut_0 = 14'b11001000100000;
9'd493   : cube_lut_0 = 14'b11001000101001;
9'd494   : cube_lut_0 = 14'b11001000110001;
9'd495   : cube_lut_0 = 14'b11001000111010;
9'd496   : cube_lut_0 = 14'b11001001000011;
9'd497   : cube_lut_0 = 14'b11001001001011;
9'd498   : cube_lut_0 = 14'b11001001010100;
9'd499   : cube_lut_0 = 14'b11001001011100;
9'd500   : cube_lut_0 = 14'b11001001100101;
9'd501   : cube_lut_0 = 14'b11001001101110;
9'd502   : cube_lut_0 = 14'b11001001110110;
9'd503   : cube_lut_0 = 14'b11001001111111;
9'd504   : cube_lut_0 = 14'b11001010000111;
9'd505   : cube_lut_0 = 14'b11001010010000;
9'd506   : cube_lut_0 = 14'b11001010011000;
9'd507   : cube_lut_0 = 14'b11001010100001;
9'd508   : cube_lut_0 = 14'b11001010101010;
9'd509   : cube_lut_0 = 14'b11001010110010;
9'd510   : cube_lut_0 = 14'b11001010111011;
9'd511   : cube_lut_0 = 14'b11001011000011;

    endcase
end

always@* begin
    
    cube_lut_1 = 0;
    
    case(i_data[8:0])
 
 9'd0   : cube_lut_1 = 14'b11001011001011;
9'd1   : cube_lut_1 = 14'b11001011010100;
9'd2   : cube_lut_1 = 14'b11001011011100;
9'd3   : cube_lut_1 = 14'b11001011100101;
9'd4   : cube_lut_1 = 14'b11001011101101;
9'd5   : cube_lut_1 = 14'b11001011110110;
9'd6   : cube_lut_1 = 14'b11001011111110;
9'd7   : cube_lut_1 = 14'b11001100000110;
9'd8   : cube_lut_1 = 14'b11001100001111;
9'd9   : cube_lut_1 = 14'b11001100010111;
9'd10   : cube_lut_1 = 14'b11001100100000;
9'd11   : cube_lut_1 = 14'b11001100101000;
9'd12   : cube_lut_1 = 14'b11001100110000;
9'd13   : cube_lut_1 = 14'b11001100111001;
9'd14   : cube_lut_1 = 14'b11001101000001;
9'd15   : cube_lut_1 = 14'b11001101001001;
9'd16   : cube_lut_1 = 14'b11001101010010;
9'd17   : cube_lut_1 = 14'b11001101011010;
9'd18   : cube_lut_1 = 14'b11001101100010;
9'd19   : cube_lut_1 = 14'b11001101101010;
9'd20   : cube_lut_1 = 14'b11001101110011;
9'd21   : cube_lut_1 = 14'b11001101111011;
9'd22   : cube_lut_1 = 14'b11001110000011;
9'd23   : cube_lut_1 = 14'b11001110001011;
9'd24   : cube_lut_1 = 14'b11001110010100;
9'd25   : cube_lut_1 = 14'b11001110011100;
9'd26   : cube_lut_1 = 14'b11001110100100;
9'd27   : cube_lut_1 = 14'b11001110101100;
9'd28   : cube_lut_1 = 14'b11001110110100;
9'd29   : cube_lut_1 = 14'b11001110111101;
9'd30   : cube_lut_1 = 14'b11001111000101;
9'd31   : cube_lut_1 = 14'b11001111001101;
9'd32   : cube_lut_1 = 14'b11001111010101;
9'd33   : cube_lut_1 = 14'b11001111011101;
9'd34   : cube_lut_1 = 14'b11001111100101;
9'd35   : cube_lut_1 = 14'b11001111101101;
9'd36   : cube_lut_1 = 14'b11001111110101;
9'd37   : cube_lut_1 = 14'b11001111111101;
9'd38   : cube_lut_1 = 14'b11010000000110;
9'd39   : cube_lut_1 = 14'b11010000001110;
9'd40   : cube_lut_1 = 14'b11010000010110;
9'd41   : cube_lut_1 = 14'b11010000011110;
9'd42   : cube_lut_1 = 14'b11010000100110;
9'd43   : cube_lut_1 = 14'b11010000101110;
9'd44   : cube_lut_1 = 14'b11010000110110;
9'd45   : cube_lut_1 = 14'b11010000111110;
9'd46   : cube_lut_1 = 14'b11010001000110;
9'd47   : cube_lut_1 = 14'b11010001001110;
9'd48   : cube_lut_1 = 14'b11010001010110;
9'd49   : cube_lut_1 = 14'b11010001011110;
9'd50   : cube_lut_1 = 14'b11010001100110;
9'd51   : cube_lut_1 = 14'b11010001101110;
9'd52   : cube_lut_1 = 14'b11010001110110;
9'd53   : cube_lut_1 = 14'b11010001111110;
9'd54   : cube_lut_1 = 14'b11010010000101;
9'd55   : cube_lut_1 = 14'b11010010001101;
9'd56   : cube_lut_1 = 14'b11010010010101;
9'd57   : cube_lut_1 = 14'b11010010011101;
9'd58   : cube_lut_1 = 14'b11010010100101;
9'd59   : cube_lut_1 = 14'b11010010101101;
9'd60   : cube_lut_1 = 14'b11010010110101;
9'd61   : cube_lut_1 = 14'b11010010111101;
9'd62   : cube_lut_1 = 14'b11010011000101;
9'd63   : cube_lut_1 = 14'b11010011001100;
9'd64   : cube_lut_1 = 14'b11010011010100;
9'd65   : cube_lut_1 = 14'b11010011011100;
9'd66   : cube_lut_1 = 14'b11010011100100;
9'd67   : cube_lut_1 = 14'b11010011101100;
9'd68   : cube_lut_1 = 14'b11010011110011;
9'd69   : cube_lut_1 = 14'b11010011111011;
9'd70   : cube_lut_1 = 14'b11010100000011;
9'd71   : cube_lut_1 = 14'b11010100001011;
9'd72   : cube_lut_1 = 14'b11010100010011;
9'd73   : cube_lut_1 = 14'b11010100011010;
9'd74   : cube_lut_1 = 14'b11010100100010;
9'd75   : cube_lut_1 = 14'b11010100101010;
9'd76   : cube_lut_1 = 14'b11010100110001;
9'd77   : cube_lut_1 = 14'b11010100111001;
9'd78   : cube_lut_1 = 14'b11010101000001;
9'd79   : cube_lut_1 = 14'b11010101001001;
9'd80   : cube_lut_1 = 14'b11010101010000;
9'd81   : cube_lut_1 = 14'b11010101011000;
9'd82   : cube_lut_1 = 14'b11010101100000;
9'd83   : cube_lut_1 = 14'b11010101100111;
9'd84   : cube_lut_1 = 14'b11010101101111;
9'd85   : cube_lut_1 = 14'b11010101110111;
9'd86   : cube_lut_1 = 14'b11010101111110;
9'd87   : cube_lut_1 = 14'b11010110000110;
9'd88   : cube_lut_1 = 14'b11010110001101;
9'd89   : cube_lut_1 = 14'b11010110010101;
9'd90   : cube_lut_1 = 14'b11010110011101;
9'd91   : cube_lut_1 = 14'b11010110100100;
9'd92   : cube_lut_1 = 14'b11010110101100;
9'd93   : cube_lut_1 = 14'b11010110110011;
9'd94   : cube_lut_1 = 14'b11010110111011;
9'd95   : cube_lut_1 = 14'b11010111000011;
9'd96   : cube_lut_1 = 14'b11010111001010;
9'd97   : cube_lut_1 = 14'b11010111010010;
9'd98   : cube_lut_1 = 14'b11010111011001;
9'd99   : cube_lut_1 = 14'b11010111100001;
9'd100   : cube_lut_1 = 14'b11010111101000;
9'd101   : cube_lut_1 = 14'b11010111110000;
9'd102   : cube_lut_1 = 14'b11010111110111;
9'd103   : cube_lut_1 = 14'b11010111111111;
9'd104   : cube_lut_1 = 14'b11011000000110;
9'd105   : cube_lut_1 = 14'b11011000001110;
9'd106   : cube_lut_1 = 14'b11011000010101;
9'd107   : cube_lut_1 = 14'b11011000011101;
9'd108   : cube_lut_1 = 14'b11011000100100;
9'd109   : cube_lut_1 = 14'b11011000101100;
9'd110   : cube_lut_1 = 14'b11011000110011;
9'd111   : cube_lut_1 = 14'b11011000111010;
9'd112   : cube_lut_1 = 14'b11011001000010;
9'd113   : cube_lut_1 = 14'b11011001001001;
9'd114   : cube_lut_1 = 14'b11011001010001;
9'd115   : cube_lut_1 = 14'b11011001011000;
9'd116   : cube_lut_1 = 14'b11011001100000;
9'd117   : cube_lut_1 = 14'b11011001100111;
9'd118   : cube_lut_1 = 14'b11011001101110;
9'd119   : cube_lut_1 = 14'b11011001110110;
9'd120   : cube_lut_1 = 14'b11011001111101;
9'd121   : cube_lut_1 = 14'b11011010000100;
9'd122   : cube_lut_1 = 14'b11011010001100;
9'd123   : cube_lut_1 = 14'b11011010010011;
9'd124   : cube_lut_1 = 14'b11011010011010;
9'd125   : cube_lut_1 = 14'b11011010100010;
9'd126   : cube_lut_1 = 14'b11011010101001;
9'd127   : cube_lut_1 = 14'b11011010110000;
9'd128   : cube_lut_1 = 14'b11011010111000;
9'd129   : cube_lut_1 = 14'b11011010111111;
9'd130   : cube_lut_1 = 14'b11011011000110;
9'd131   : cube_lut_1 = 14'b11011011001101;
9'd132   : cube_lut_1 = 14'b11011011010101;
9'd133   : cube_lut_1 = 14'b11011011011100;
9'd134   : cube_lut_1 = 14'b11011011100011;
9'd135   : cube_lut_1 = 14'b11011011101011;
9'd136   : cube_lut_1 = 14'b11011011110010;
9'd137   : cube_lut_1 = 14'b11011011111001;
9'd138   : cube_lut_1 = 14'b11011100000000;
9'd139   : cube_lut_1 = 14'b11011100000111;
9'd140   : cube_lut_1 = 14'b11011100001111;
9'd141   : cube_lut_1 = 14'b11011100010110;
9'd142   : cube_lut_1 = 14'b11011100011101;
9'd143   : cube_lut_1 = 14'b11011100100100;
9'd144   : cube_lut_1 = 14'b11011100101011;
9'd145   : cube_lut_1 = 14'b11011100110011;
9'd146   : cube_lut_1 = 14'b11011100111010;
9'd147   : cube_lut_1 = 14'b11011101000001;
9'd148   : cube_lut_1 = 14'b11011101001000;
9'd149   : cube_lut_1 = 14'b11011101001111;
9'd150   : cube_lut_1 = 14'b11011101010110;
9'd151   : cube_lut_1 = 14'b11011101011101;
9'd152   : cube_lut_1 = 14'b11011101100101;
9'd153   : cube_lut_1 = 14'b11011101101100;
9'd154   : cube_lut_1 = 14'b11011101110011;
9'd155   : cube_lut_1 = 14'b11011101111010;
9'd156   : cube_lut_1 = 14'b11011110000001;
9'd157   : cube_lut_1 = 14'b11011110001000;
9'd158   : cube_lut_1 = 14'b11011110001111;
9'd159   : cube_lut_1 = 14'b11011110010110;
9'd160   : cube_lut_1 = 14'b11011110011101;
9'd161   : cube_lut_1 = 14'b11011110100100;
9'd162   : cube_lut_1 = 14'b11011110101011;
9'd163   : cube_lut_1 = 14'b11011110110010;
9'd164   : cube_lut_1 = 14'b11011110111001;
9'd165   : cube_lut_1 = 14'b11011111000001;
9'd166   : cube_lut_1 = 14'b11011111001000;
9'd167   : cube_lut_1 = 14'b11011111001111;
9'd168   : cube_lut_1 = 14'b11011111010110;
9'd169   : cube_lut_1 = 14'b11011111011101;
9'd170   : cube_lut_1 = 14'b11011111100100;
9'd171   : cube_lut_1 = 14'b11011111101011;
9'd172   : cube_lut_1 = 14'b11011111110010;
9'd173   : cube_lut_1 = 14'b11011111111001;
9'd174   : cube_lut_1 = 14'b11100000000000;
9'd175   : cube_lut_1 = 14'b11100000000110;
9'd176   : cube_lut_1 = 14'b11100000001101;
9'd177   : cube_lut_1 = 14'b11100000010100;
9'd178   : cube_lut_1 = 14'b11100000011011;
9'd179   : cube_lut_1 = 14'b11100000100010;
9'd180   : cube_lut_1 = 14'b11100000101001;
9'd181   : cube_lut_1 = 14'b11100000110000;
9'd182   : cube_lut_1 = 14'b11100000110111;
9'd183   : cube_lut_1 = 14'b11100000111110;
9'd184   : cube_lut_1 = 14'b11100001000101;
9'd185   : cube_lut_1 = 14'b11100001001100;
9'd186   : cube_lut_1 = 14'b11100001010011;
9'd187   : cube_lut_1 = 14'b11100001011001;
9'd188   : cube_lut_1 = 14'b11100001100000;
9'd189   : cube_lut_1 = 14'b11100001100111;
9'd190   : cube_lut_1 = 14'b11100001101110;
9'd191   : cube_lut_1 = 14'b11100001110101;
9'd192   : cube_lut_1 = 14'b11100001111100;
9'd193   : cube_lut_1 = 14'b11100010000011;
9'd194   : cube_lut_1 = 14'b11100010001001;
9'd195   : cube_lut_1 = 14'b11100010010000;
9'd196   : cube_lut_1 = 14'b11100010010111;
9'd197   : cube_lut_1 = 14'b11100010011110;
9'd198   : cube_lut_1 = 14'b11100010100101;
9'd199   : cube_lut_1 = 14'b11100010101100;
9'd200   : cube_lut_1 = 14'b11100010110010;
9'd201   : cube_lut_1 = 14'b11100010111001;
9'd202   : cube_lut_1 = 14'b11100011000000;
9'd203   : cube_lut_1 = 14'b11100011000111;
9'd204   : cube_lut_1 = 14'b11100011001110;
9'd205   : cube_lut_1 = 14'b11100011010100;
9'd206   : cube_lut_1 = 14'b11100011011011;
9'd207   : cube_lut_1 = 14'b11100011100010;
9'd208   : cube_lut_1 = 14'b11100011101001;
9'd209   : cube_lut_1 = 14'b11100011101111;
9'd210   : cube_lut_1 = 14'b11100011110110;
9'd211   : cube_lut_1 = 14'b11100011111101;
9'd212   : cube_lut_1 = 14'b11100100000011;
9'd213   : cube_lut_1 = 14'b11100100001010;
9'd214   : cube_lut_1 = 14'b11100100010001;
9'd215   : cube_lut_1 = 14'b11100100011000;
9'd216   : cube_lut_1 = 14'b11100100011110;
9'd217   : cube_lut_1 = 14'b11100100100101;
9'd218   : cube_lut_1 = 14'b11100100101100;
9'd219   : cube_lut_1 = 14'b11100100110010;
9'd220   : cube_lut_1 = 14'b11100100111001;
9'd221   : cube_lut_1 = 14'b11100101000000;
9'd222   : cube_lut_1 = 14'b11100101000110;
9'd223   : cube_lut_1 = 14'b11100101001101;
9'd224   : cube_lut_1 = 14'b11100101010100;
9'd225   : cube_lut_1 = 14'b11100101011010;
9'd226   : cube_lut_1 = 14'b11100101100001;
9'd227   : cube_lut_1 = 14'b11100101101000;
9'd228   : cube_lut_1 = 14'b11100101101110;
9'd229   : cube_lut_1 = 14'b11100101110101;
9'd230   : cube_lut_1 = 14'b11100101111011;
9'd231   : cube_lut_1 = 14'b11100110000010;
9'd232   : cube_lut_1 = 14'b11100110001001;
9'd233   : cube_lut_1 = 14'b11100110001111;
9'd234   : cube_lut_1 = 14'b11100110010110;
9'd235   : cube_lut_1 = 14'b11100110011100;
9'd236   : cube_lut_1 = 14'b11100110100011;
9'd237   : cube_lut_1 = 14'b11100110101010;
9'd238   : cube_lut_1 = 14'b11100110110000;
9'd239   : cube_lut_1 = 14'b11100110110111;
9'd240   : cube_lut_1 = 14'b11100110111101;
9'd241   : cube_lut_1 = 14'b11100111000100;
9'd242   : cube_lut_1 = 14'b11100111001010;
9'd243   : cube_lut_1 = 14'b11100111010001;
9'd244   : cube_lut_1 = 14'b11100111010111;
9'd245   : cube_lut_1 = 14'b11100111011110;
9'd246   : cube_lut_1 = 14'b11100111100100;
9'd247   : cube_lut_1 = 14'b11100111101011;
9'd248   : cube_lut_1 = 14'b11100111110001;
9'd249   : cube_lut_1 = 14'b11100111111000;
9'd250   : cube_lut_1 = 14'b11100111111110;
9'd251   : cube_lut_1 = 14'b11101000000101;
9'd252   : cube_lut_1 = 14'b11101000001011;
9'd253   : cube_lut_1 = 14'b11101000010010;
9'd254   : cube_lut_1 = 14'b11101000011000;
9'd255   : cube_lut_1 = 14'b11101000011111;
9'd256   : cube_lut_1 = 14'b11101000100101;
9'd257   : cube_lut_1 = 14'b11101000101100;
9'd258   : cube_lut_1 = 14'b11101000110010;
9'd259   : cube_lut_1 = 14'b11101000111001;
9'd260   : cube_lut_1 = 14'b11101000111111;
9'd261   : cube_lut_1 = 14'b11101001000110;
9'd262   : cube_lut_1 = 14'b11101001001100;
9'd263   : cube_lut_1 = 14'b11101001010010;
9'd264   : cube_lut_1 = 14'b11101001011001;
9'd265   : cube_lut_1 = 14'b11101001011111;
9'd266   : cube_lut_1 = 14'b11101001100110;
9'd267   : cube_lut_1 = 14'b11101001101100;
9'd268   : cube_lut_1 = 14'b11101001110010;
9'd269   : cube_lut_1 = 14'b11101001111001;
9'd270   : cube_lut_1 = 14'b11101001111111;
9'd271   : cube_lut_1 = 14'b11101010000110;
9'd272   : cube_lut_1 = 14'b11101010001100;
9'd273   : cube_lut_1 = 14'b11101010010010;
9'd274   : cube_lut_1 = 14'b11101010011001;
9'd275   : cube_lut_1 = 14'b11101010011111;
9'd276   : cube_lut_1 = 14'b11101010100101;
9'd277   : cube_lut_1 = 14'b11101010101100;
9'd278   : cube_lut_1 = 14'b11101010110010;
9'd279   : cube_lut_1 = 14'b11101010111000;
9'd280   : cube_lut_1 = 14'b11101010111111;
9'd281   : cube_lut_1 = 14'b11101011000101;
9'd282   : cube_lut_1 = 14'b11101011001011;
9'd283   : cube_lut_1 = 14'b11101011010010;
9'd284   : cube_lut_1 = 14'b11101011011000;
9'd285   : cube_lut_1 = 14'b11101011011110;
9'd286   : cube_lut_1 = 14'b11101011100101;
9'd287   : cube_lut_1 = 14'b11101011101011;
9'd288   : cube_lut_1 = 14'b11101011110001;
9'd289   : cube_lut_1 = 14'b11101011111000;
9'd290   : cube_lut_1 = 14'b11101011111110;
9'd291   : cube_lut_1 = 14'b11101100000100;
9'd292   : cube_lut_1 = 14'b11101100001010;
9'd293   : cube_lut_1 = 14'b11101100010001;
9'd294   : cube_lut_1 = 14'b11101100010111;
9'd295   : cube_lut_1 = 14'b11101100011101;
9'd296   : cube_lut_1 = 14'b11101100100011;
9'd297   : cube_lut_1 = 14'b11101100101010;
9'd298   : cube_lut_1 = 14'b11101100110000;
9'd299   : cube_lut_1 = 14'b11101100110110;
9'd300   : cube_lut_1 = 14'b11101100111100;
9'd301   : cube_lut_1 = 14'b11101101000011;
9'd302   : cube_lut_1 = 14'b11101101001001;
9'd303   : cube_lut_1 = 14'b11101101001111;
9'd304   : cube_lut_1 = 14'b11101101010101;
9'd305   : cube_lut_1 = 14'b11101101011011;
9'd306   : cube_lut_1 = 14'b11101101100010;
9'd307   : cube_lut_1 = 14'b11101101101000;
9'd308   : cube_lut_1 = 14'b11101101101110;
9'd309   : cube_lut_1 = 14'b11101101110100;
9'd310   : cube_lut_1 = 14'b11101101111010;
9'd311   : cube_lut_1 = 14'b11101110000001;
9'd312   : cube_lut_1 = 14'b11101110000111;
9'd313   : cube_lut_1 = 14'b11101110001101;
9'd314   : cube_lut_1 = 14'b11101110010011;
9'd315   : cube_lut_1 = 14'b11101110011001;
9'd316   : cube_lut_1 = 14'b11101110011111;
9'd317   : cube_lut_1 = 14'b11101110100101;
9'd318   : cube_lut_1 = 14'b11101110101100;
9'd319   : cube_lut_1 = 14'b11101110110010;
9'd320   : cube_lut_1 = 14'b11101110111000;
9'd321   : cube_lut_1 = 14'b11101110111110;
9'd322   : cube_lut_1 = 14'b11101111000100;
9'd323   : cube_lut_1 = 14'b11101111001010;
9'd324   : cube_lut_1 = 14'b11101111010000;
9'd325   : cube_lut_1 = 14'b11101111010110;
9'd326   : cube_lut_1 = 14'b11101111011101;
9'd327   : cube_lut_1 = 14'b11101111100011;
9'd328   : cube_lut_1 = 14'b11101111101001;
9'd329   : cube_lut_1 = 14'b11101111101111;
9'd330   : cube_lut_1 = 14'b11101111110101;
9'd331   : cube_lut_1 = 14'b11101111111011;
9'd332   : cube_lut_1 = 14'b11110000000001;
9'd333   : cube_lut_1 = 14'b11110000000111;
9'd334   : cube_lut_1 = 14'b11110000001101;
9'd335   : cube_lut_1 = 14'b11110000010011;
9'd336   : cube_lut_1 = 14'b11110000011001;
9'd337   : cube_lut_1 = 14'b11110000011111;
9'd338   : cube_lut_1 = 14'b11110000100101;
9'd339   : cube_lut_1 = 14'b11110000101011;
9'd340   : cube_lut_1 = 14'b11110000110001;
9'd341   : cube_lut_1 = 14'b11110000110111;
9'd342   : cube_lut_1 = 14'b11110000111101;
9'd343   : cube_lut_1 = 14'b11110001000011;
9'd344   : cube_lut_1 = 14'b11110001001001;
9'd345   : cube_lut_1 = 14'b11110001001111;
9'd346   : cube_lut_1 = 14'b11110001010101;
9'd347   : cube_lut_1 = 14'b11110001011011;
9'd348   : cube_lut_1 = 14'b11110001100001;
9'd349   : cube_lut_1 = 14'b11110001100111;
9'd350   : cube_lut_1 = 14'b11110001101101;
9'd351   : cube_lut_1 = 14'b11110001110011;
9'd352   : cube_lut_1 = 14'b11110001111001;
9'd353   : cube_lut_1 = 14'b11110001111111;
9'd354   : cube_lut_1 = 14'b11110010000101;
9'd355   : cube_lut_1 = 14'b11110010001011;
9'd356   : cube_lut_1 = 14'b11110010010001;
9'd357   : cube_lut_1 = 14'b11110010010111;
9'd358   : cube_lut_1 = 14'b11110010011101;
9'd359   : cube_lut_1 = 14'b11110010100011;
9'd360   : cube_lut_1 = 14'b11110010101001;
9'd361   : cube_lut_1 = 14'b11110010101111;
9'd362   : cube_lut_1 = 14'b11110010110101;
9'd363   : cube_lut_1 = 14'b11110010111011;
9'd364   : cube_lut_1 = 14'b11110011000001;
9'd365   : cube_lut_1 = 14'b11110011000111;
9'd366   : cube_lut_1 = 14'b11110011001101;
9'd367   : cube_lut_1 = 14'b11110011010010;
9'd368   : cube_lut_1 = 14'b11110011011000;
9'd369   : cube_lut_1 = 14'b11110011011110;
9'd370   : cube_lut_1 = 14'b11110011100100;
9'd371   : cube_lut_1 = 14'b11110011101010;
9'd372   : cube_lut_1 = 14'b11110011110000;
9'd373   : cube_lut_1 = 14'b11110011110110;
9'd374   : cube_lut_1 = 14'b11110011111100;
9'd375   : cube_lut_1 = 14'b11110100000010;
9'd376   : cube_lut_1 = 14'b11110100000111;
9'd377   : cube_lut_1 = 14'b11110100001101;
9'd378   : cube_lut_1 = 14'b11110100010011;
9'd379   : cube_lut_1 = 14'b11110100011001;
9'd380   : cube_lut_1 = 14'b11110100011111;
9'd381   : cube_lut_1 = 14'b11110100100101;
9'd382   : cube_lut_1 = 14'b11110100101011;
9'd383   : cube_lut_1 = 14'b11110100110000;
9'd384   : cube_lut_1 = 14'b11110100110110;
9'd385   : cube_lut_1 = 14'b11110100111100;
9'd386   : cube_lut_1 = 14'b11110101000010;
9'd387   : cube_lut_1 = 14'b11110101001000;
9'd388   : cube_lut_1 = 14'b11110101001110;
9'd389   : cube_lut_1 = 14'b11110101010011;
9'd390   : cube_lut_1 = 14'b11110101011001;
9'd391   : cube_lut_1 = 14'b11110101011111;
9'd392   : cube_lut_1 = 14'b11110101100101;
9'd393   : cube_lut_1 = 14'b11110101101011;
9'd394   : cube_lut_1 = 14'b11110101110000;
9'd395   : cube_lut_1 = 14'b11110101110110;
9'd396   : cube_lut_1 = 14'b11110101111100;
9'd397   : cube_lut_1 = 14'b11110110000010;
9'd398   : cube_lut_1 = 14'b11110110000111;
9'd399   : cube_lut_1 = 14'b11110110001101;
9'd400   : cube_lut_1 = 14'b11110110010011;
9'd401   : cube_lut_1 = 14'b11110110011001;
9'd402   : cube_lut_1 = 14'b11110110011110;
9'd403   : cube_lut_1 = 14'b11110110100100;
9'd404   : cube_lut_1 = 14'b11110110101010;
9'd405   : cube_lut_1 = 14'b11110110110000;
9'd406   : cube_lut_1 = 14'b11110110110101;
9'd407   : cube_lut_1 = 14'b11110110111011;
9'd408   : cube_lut_1 = 14'b11110111000001;
9'd409   : cube_lut_1 = 14'b11110111000111;
9'd410   : cube_lut_1 = 14'b11110111001100;
9'd411   : cube_lut_1 = 14'b11110111010010;
9'd412   : cube_lut_1 = 14'b11110111011000;
9'd413   : cube_lut_1 = 14'b11110111011110;
9'd414   : cube_lut_1 = 14'b11110111100011;
9'd415   : cube_lut_1 = 14'b11110111101001;
9'd416   : cube_lut_1 = 14'b11110111101111;
9'd417   : cube_lut_1 = 14'b11110111110100;
9'd418   : cube_lut_1 = 14'b11110111111010;
9'd419   : cube_lut_1 = 14'b11111000000000;
9'd420   : cube_lut_1 = 14'b11111000000101;
9'd421   : cube_lut_1 = 14'b11111000001011;
9'd422   : cube_lut_1 = 14'b11111000010001;
9'd423   : cube_lut_1 = 14'b11111000010110;
9'd424   : cube_lut_1 = 14'b11111000011100;
9'd425   : cube_lut_1 = 14'b11111000100010;
9'd426   : cube_lut_1 = 14'b11111000100111;
9'd427   : cube_lut_1 = 14'b11111000101101;
9'd428   : cube_lut_1 = 14'b11111000110011;
9'd429   : cube_lut_1 = 14'b11111000111000;
9'd430   : cube_lut_1 = 14'b11111000111110;
9'd431   : cube_lut_1 = 14'b11111001000100;
9'd432   : cube_lut_1 = 14'b11111001001001;
9'd433   : cube_lut_1 = 14'b11111001001111;
9'd434   : cube_lut_1 = 14'b11111001010100;
9'd435   : cube_lut_1 = 14'b11111001011010;
9'd436   : cube_lut_1 = 14'b11111001100000;
9'd437   : cube_lut_1 = 14'b11111001100101;
9'd438   : cube_lut_1 = 14'b11111001101011;
9'd439   : cube_lut_1 = 14'b11111001110001;
9'd440   : cube_lut_1 = 14'b11111001110110;
9'd441   : cube_lut_1 = 14'b11111001111100;
9'd442   : cube_lut_1 = 14'b11111010000001;
9'd443   : cube_lut_1 = 14'b11111010000111;
9'd444   : cube_lut_1 = 14'b11111010001100;
9'd445   : cube_lut_1 = 14'b11111010010010;
9'd446   : cube_lut_1 = 14'b11111010011000;
9'd447   : cube_lut_1 = 14'b11111010011101;
9'd448   : cube_lut_1 = 14'b11111010100011;
9'd449   : cube_lut_1 = 14'b11111010101000;
9'd450   : cube_lut_1 = 14'b11111010101110;
9'd451   : cube_lut_1 = 14'b11111010110011;
9'd452   : cube_lut_1 = 14'b11111010111001;
9'd453   : cube_lut_1 = 14'b11111010111111;
9'd454   : cube_lut_1 = 14'b11111011000100;
9'd455   : cube_lut_1 = 14'b11111011001010;
9'd456   : cube_lut_1 = 14'b11111011001111;
9'd457   : cube_lut_1 = 14'b11111011010101;
9'd458   : cube_lut_1 = 14'b11111011011010;
9'd459   : cube_lut_1 = 14'b11111011100000;
9'd460   : cube_lut_1 = 14'b11111011100101;
9'd461   : cube_lut_1 = 14'b11111011101011;
9'd462   : cube_lut_1 = 14'b11111011110000;
9'd463   : cube_lut_1 = 14'b11111011110110;
9'd464   : cube_lut_1 = 14'b11111011111011;
9'd465   : cube_lut_1 = 14'b11111100000001;
9'd466   : cube_lut_1 = 14'b11111100000110;
9'd467   : cube_lut_1 = 14'b11111100001100;
9'd468   : cube_lut_1 = 14'b11111100010001;
9'd469   : cube_lut_1 = 14'b11111100010111;
9'd470   : cube_lut_1 = 14'b11111100011100;
9'd471   : cube_lut_1 = 14'b11111100100010;
9'd472   : cube_lut_1 = 14'b11111100100111;
9'd473   : cube_lut_1 = 14'b11111100101101;
9'd474   : cube_lut_1 = 14'b11111100110010;
9'd475   : cube_lut_1 = 14'b11111100111000;
9'd476   : cube_lut_1 = 14'b11111100111101;
9'd477   : cube_lut_1 = 14'b11111101000011;
9'd478   : cube_lut_1 = 14'b11111101001000;
9'd479   : cube_lut_1 = 14'b11111101001110;
9'd480   : cube_lut_1 = 14'b11111101010011;
9'd481   : cube_lut_1 = 14'b11111101011000;
9'd482   : cube_lut_1 = 14'b11111101011110;
9'd483   : cube_lut_1 = 14'b11111101100011;
9'd484   : cube_lut_1 = 14'b11111101101001;
9'd485   : cube_lut_1 = 14'b11111101101110;
9'd486   : cube_lut_1 = 14'b11111101110100;
9'd487   : cube_lut_1 = 14'b11111101111001;
9'd488   : cube_lut_1 = 14'b11111101111110;
9'd489   : cube_lut_1 = 14'b11111110000100;
9'd490   : cube_lut_1 = 14'b11111110001001;
9'd491   : cube_lut_1 = 14'b11111110001111;
9'd492   : cube_lut_1 = 14'b11111110010100;
9'd493   : cube_lut_1 = 14'b11111110011010;
9'd494   : cube_lut_1 = 14'b11111110011111;
9'd495   : cube_lut_1 = 14'b11111110100100;
9'd496   : cube_lut_1 = 14'b11111110101010;
9'd497   : cube_lut_1 = 14'b11111110101111;
9'd498   : cube_lut_1 = 14'b11111110110100;
9'd499   : cube_lut_1 = 14'b11111110111010;
9'd500   : cube_lut_1 = 14'b11111110111111;
9'd501   : cube_lut_1 = 14'b11111111000101;
9'd502   : cube_lut_1 = 14'b11111111001010;
9'd503   : cube_lut_1 = 14'b11111111001111;
9'd504   : cube_lut_1 = 14'b11111111010101;
9'd505   : cube_lut_1 = 14'b11111111011010;
9'd506   : cube_lut_1 = 14'b11111111011111;
9'd507   : cube_lut_1 = 14'b11111111100101;
9'd508   : cube_lut_1 = 14'b11111111101010;
9'd509   : cube_lut_1 = 14'b11111111101111;
9'd510   : cube_lut_1 = 14'b11111111110101;
9'd511   : cube_lut_1 = 14'b11111111111010;

    endcase
end

always@* begin
    
    cube_lut_2 = 0;
    
    case(i_data[8:0])
 
 9'd0   : cube_lut_2 = 14'b10000000000000;
9'd1   : cube_lut_2 = 14'b10000000000010;
9'd2   : cube_lut_2 = 14'b10000000000101;
9'd3   : cube_lut_2 = 14'b10000000000111;
9'd4   : cube_lut_2 = 14'b10000000001010;
9'd5   : cube_lut_2 = 14'b10000000001101;
9'd6   : cube_lut_2 = 14'b10000000001111;
9'd7   : cube_lut_2 = 14'b10000000010010;
9'd8   : cube_lut_2 = 14'b10000000010101;
9'd9   : cube_lut_2 = 14'b10000000010111;
9'd10   : cube_lut_2 = 14'b10000000011010;
9'd11   : cube_lut_2 = 14'b10000000011101;
9'd12   : cube_lut_2 = 14'b10000000011111;
9'd13   : cube_lut_2 = 14'b10000000100010;
9'd14   : cube_lut_2 = 14'b10000000100101;
9'd15   : cube_lut_2 = 14'b10000000100111;
9'd16   : cube_lut_2 = 14'b10000000101010;
9'd17   : cube_lut_2 = 14'b10000000101101;
9'd18   : cube_lut_2 = 14'b10000000101111;
9'd19   : cube_lut_2 = 14'b10000000110010;
9'd20   : cube_lut_2 = 14'b10000000110100;
9'd21   : cube_lut_2 = 14'b10000000110111;
9'd22   : cube_lut_2 = 14'b10000000111010;
9'd23   : cube_lut_2 = 14'b10000000111100;
9'd24   : cube_lut_2 = 14'b10000000111111;
9'd25   : cube_lut_2 = 14'b10000001000010;
9'd26   : cube_lut_2 = 14'b10000001000100;
9'd27   : cube_lut_2 = 14'b10000001000111;
9'd28   : cube_lut_2 = 14'b10000001001001;
9'd29   : cube_lut_2 = 14'b10000001001100;
9'd30   : cube_lut_2 = 14'b10000001001111;
9'd31   : cube_lut_2 = 14'b10000001010001;
9'd32   : cube_lut_2 = 14'b10000001010100;
9'd33   : cube_lut_2 = 14'b10000001010111;
9'd34   : cube_lut_2 = 14'b10000001011001;
9'd35   : cube_lut_2 = 14'b10000001011100;
9'd36   : cube_lut_2 = 14'b10000001011110;
9'd37   : cube_lut_2 = 14'b10000001100001;
9'd38   : cube_lut_2 = 14'b10000001100100;
9'd39   : cube_lut_2 = 14'b10000001100110;
9'd40   : cube_lut_2 = 14'b10000001101001;
9'd41   : cube_lut_2 = 14'b10000001101011;
9'd42   : cube_lut_2 = 14'b10000001101110;
9'd43   : cube_lut_2 = 14'b10000001110001;
9'd44   : cube_lut_2 = 14'b10000001110011;
9'd45   : cube_lut_2 = 14'b10000001110110;
9'd46   : cube_lut_2 = 14'b10000001111000;
9'd47   : cube_lut_2 = 14'b10000001111011;
9'd48   : cube_lut_2 = 14'b10000001111110;
9'd49   : cube_lut_2 = 14'b10000010000000;
9'd50   : cube_lut_2 = 14'b10000010000011;
9'd51   : cube_lut_2 = 14'b10000010000101;
9'd52   : cube_lut_2 = 14'b10000010001000;
9'd53   : cube_lut_2 = 14'b10000010001010;
9'd54   : cube_lut_2 = 14'b10000010001101;
9'd55   : cube_lut_2 = 14'b10000010010000;
9'd56   : cube_lut_2 = 14'b10000010010010;
9'd57   : cube_lut_2 = 14'b10000010010101;
9'd58   : cube_lut_2 = 14'b10000010010111;
9'd59   : cube_lut_2 = 14'b10000010011010;
9'd60   : cube_lut_2 = 14'b10000010011100;
9'd61   : cube_lut_2 = 14'b10000010011111;
9'd62   : cube_lut_2 = 14'b10000010100010;
9'd63   : cube_lut_2 = 14'b10000010100100;
9'd64   : cube_lut_2 = 14'b10000010100111;
9'd65   : cube_lut_2 = 14'b10000010101001;
9'd66   : cube_lut_2 = 14'b10000010101100;
9'd67   : cube_lut_2 = 14'b10000010101110;
9'd68   : cube_lut_2 = 14'b10000010110001;
9'd69   : cube_lut_2 = 14'b10000010110100;
9'd70   : cube_lut_2 = 14'b10000010110110;
9'd71   : cube_lut_2 = 14'b10000010111001;
9'd72   : cube_lut_2 = 14'b10000010111011;
9'd73   : cube_lut_2 = 14'b10000010111110;
9'd74   : cube_lut_2 = 14'b10000011000000;
9'd75   : cube_lut_2 = 14'b10000011000011;
9'd76   : cube_lut_2 = 14'b10000011000101;
9'd77   : cube_lut_2 = 14'b10000011001000;
9'd78   : cube_lut_2 = 14'b10000011001010;
9'd79   : cube_lut_2 = 14'b10000011001101;
9'd80   : cube_lut_2 = 14'b10000011010000;
9'd81   : cube_lut_2 = 14'b10000011010010;
9'd82   : cube_lut_2 = 14'b10000011010101;
9'd83   : cube_lut_2 = 14'b10000011010111;
9'd84   : cube_lut_2 = 14'b10000011011010;
9'd85   : cube_lut_2 = 14'b10000011011100;
9'd86   : cube_lut_2 = 14'b10000011011111;
9'd87   : cube_lut_2 = 14'b10000011100001;
9'd88   : cube_lut_2 = 14'b10000011100100;
9'd89   : cube_lut_2 = 14'b10000011100110;
9'd90   : cube_lut_2 = 14'b10000011101001;
9'd91   : cube_lut_2 = 14'b10000011101011;
9'd92   : cube_lut_2 = 14'b10000011101110;
9'd93   : cube_lut_2 = 14'b10000011110000;
9'd94   : cube_lut_2 = 14'b10000011110011;
9'd95   : cube_lut_2 = 14'b10000011110101;
9'd96   : cube_lut_2 = 14'b10000011111000;
9'd97   : cube_lut_2 = 14'b10000011111010;
9'd98   : cube_lut_2 = 14'b10000011111101;
9'd99   : cube_lut_2 = 14'b10000011111111;
9'd100   : cube_lut_2 = 14'b10000100000010;
9'd101   : cube_lut_2 = 14'b10000100000100;
9'd102   : cube_lut_2 = 14'b10000100000111;
9'd103   : cube_lut_2 = 14'b10000100001001;
9'd104   : cube_lut_2 = 14'b10000100001100;
9'd105   : cube_lut_2 = 14'b10000100001110;
9'd106   : cube_lut_2 = 14'b10000100010001;
9'd107   : cube_lut_2 = 14'b10000100010011;
9'd108   : cube_lut_2 = 14'b10000100010110;
9'd109   : cube_lut_2 = 14'b10000100011000;
9'd110   : cube_lut_2 = 14'b10000100011011;
9'd111   : cube_lut_2 = 14'b10000100011101;
9'd112   : cube_lut_2 = 14'b10000100100000;
9'd113   : cube_lut_2 = 14'b10000100100010;
9'd114   : cube_lut_2 = 14'b10000100100101;
9'd115   : cube_lut_2 = 14'b10000100100111;
9'd116   : cube_lut_2 = 14'b10000100101010;
9'd117   : cube_lut_2 = 14'b10000100101100;
9'd118   : cube_lut_2 = 14'b10000100101111;
9'd119   : cube_lut_2 = 14'b10000100110001;
9'd120   : cube_lut_2 = 14'b10000100110100;
9'd121   : cube_lut_2 = 14'b10000100110110;
9'd122   : cube_lut_2 = 14'b10000100111001;
9'd123   : cube_lut_2 = 14'b10000100111011;
9'd124   : cube_lut_2 = 14'b10000100111110;
9'd125   : cube_lut_2 = 14'b10000101000000;
9'd126   : cube_lut_2 = 14'b10000101000011;
9'd127   : cube_lut_2 = 14'b10000101000101;
9'd128   : cube_lut_2 = 14'b10000101001000;
9'd129   : cube_lut_2 = 14'b10000101001010;
9'd130   : cube_lut_2 = 14'b10000101001100;
9'd131   : cube_lut_2 = 14'b10000101001111;
9'd132   : cube_lut_2 = 14'b10000101010001;
9'd133   : cube_lut_2 = 14'b10000101010100;
9'd134   : cube_lut_2 = 14'b10000101010110;
9'd135   : cube_lut_2 = 14'b10000101011001;
9'd136   : cube_lut_2 = 14'b10000101011011;
9'd137   : cube_lut_2 = 14'b10000101011110;
9'd138   : cube_lut_2 = 14'b10000101100000;
9'd139   : cube_lut_2 = 14'b10000101100011;
9'd140   : cube_lut_2 = 14'b10000101100101;
9'd141   : cube_lut_2 = 14'b10000101100111;
9'd142   : cube_lut_2 = 14'b10000101101010;
9'd143   : cube_lut_2 = 14'b10000101101100;
9'd144   : cube_lut_2 = 14'b10000101101111;
9'd145   : cube_lut_2 = 14'b10000101110001;
9'd146   : cube_lut_2 = 14'b10000101110100;
9'd147   : cube_lut_2 = 14'b10000101110110;
9'd148   : cube_lut_2 = 14'b10000101111001;
9'd149   : cube_lut_2 = 14'b10000101111011;
9'd150   : cube_lut_2 = 14'b10000101111101;
9'd151   : cube_lut_2 = 14'b10000110000000;
9'd152   : cube_lut_2 = 14'b10000110000010;
9'd153   : cube_lut_2 = 14'b10000110000101;
9'd154   : cube_lut_2 = 14'b10000110000111;
9'd155   : cube_lut_2 = 14'b10000110001010;
9'd156   : cube_lut_2 = 14'b10000110001100;
9'd157   : cube_lut_2 = 14'b10000110001110;
9'd158   : cube_lut_2 = 14'b10000110010001;
9'd159   : cube_lut_2 = 14'b10000110010011;
9'd160   : cube_lut_2 = 14'b10000110010110;
9'd161   : cube_lut_2 = 14'b10000110011000;
9'd162   : cube_lut_2 = 14'b10000110011011;
9'd163   : cube_lut_2 = 14'b10000110011101;
9'd164   : cube_lut_2 = 14'b10000110011111;
9'd165   : cube_lut_2 = 14'b10000110100010;
9'd166   : cube_lut_2 = 14'b10000110100100;
9'd167   : cube_lut_2 = 14'b10000110100111;
9'd168   : cube_lut_2 = 14'b10000110101001;
9'd169   : cube_lut_2 = 14'b10000110101011;
9'd170   : cube_lut_2 = 14'b10000110101110;
9'd171   : cube_lut_2 = 14'b10000110110000;
9'd172   : cube_lut_2 = 14'b10000110110011;
9'd173   : cube_lut_2 = 14'b10000110110101;
9'd174   : cube_lut_2 = 14'b10000110110111;
9'd175   : cube_lut_2 = 14'b10000110111010;
9'd176   : cube_lut_2 = 14'b10000110111100;
9'd177   : cube_lut_2 = 14'b10000110111111;
9'd178   : cube_lut_2 = 14'b10000111000001;
9'd179   : cube_lut_2 = 14'b10000111000011;
9'd180   : cube_lut_2 = 14'b10000111000110;
9'd181   : cube_lut_2 = 14'b10000111001000;
9'd182   : cube_lut_2 = 14'b10000111001011;
9'd183   : cube_lut_2 = 14'b10000111001101;
9'd184   : cube_lut_2 = 14'b10000111001111;
9'd185   : cube_lut_2 = 14'b10000111010010;
9'd186   : cube_lut_2 = 14'b10000111010100;
9'd187   : cube_lut_2 = 14'b10000111010111;
9'd188   : cube_lut_2 = 14'b10000111011001;
9'd189   : cube_lut_2 = 14'b10000111011011;
9'd190   : cube_lut_2 = 14'b10000111011110;
9'd191   : cube_lut_2 = 14'b10000111100000;
9'd192   : cube_lut_2 = 14'b10000111100010;
9'd193   : cube_lut_2 = 14'b10000111100101;
9'd194   : cube_lut_2 = 14'b10000111100111;
9'd195   : cube_lut_2 = 14'b10000111101010;
9'd196   : cube_lut_2 = 14'b10000111101100;
9'd197   : cube_lut_2 = 14'b10000111101110;
9'd198   : cube_lut_2 = 14'b10000111110001;
9'd199   : cube_lut_2 = 14'b10000111110011;
9'd200   : cube_lut_2 = 14'b10000111110101;
9'd201   : cube_lut_2 = 14'b10000111111000;
9'd202   : cube_lut_2 = 14'b10000111111010;
9'd203   : cube_lut_2 = 14'b10000111111101;
9'd204   : cube_lut_2 = 14'b10000111111111;
9'd205   : cube_lut_2 = 14'b10001000000001;
9'd206   : cube_lut_2 = 14'b10001000000100;
9'd207   : cube_lut_2 = 14'b10001000000110;
9'd208   : cube_lut_2 = 14'b10001000001000;
9'd209   : cube_lut_2 = 14'b10001000001011;
9'd210   : cube_lut_2 = 14'b10001000001101;
9'd211   : cube_lut_2 = 14'b10001000001111;
9'd212   : cube_lut_2 = 14'b10001000010010;
9'd213   : cube_lut_2 = 14'b10001000010100;
9'd214   : cube_lut_2 = 14'b10001000010110;
9'd215   : cube_lut_2 = 14'b10001000011001;
9'd216   : cube_lut_2 = 14'b10001000011011;
9'd217   : cube_lut_2 = 14'b10001000011110;
9'd218   : cube_lut_2 = 14'b10001000100000;
9'd219   : cube_lut_2 = 14'b10001000100010;
9'd220   : cube_lut_2 = 14'b10001000100101;
9'd221   : cube_lut_2 = 14'b10001000100111;
9'd222   : cube_lut_2 = 14'b10001000101001;
9'd223   : cube_lut_2 = 14'b10001000101100;
9'd224   : cube_lut_2 = 14'b10001000101110;
9'd225   : cube_lut_2 = 14'b10001000110000;
9'd226   : cube_lut_2 = 14'b10001000110011;
9'd227   : cube_lut_2 = 14'b10001000110101;
9'd228   : cube_lut_2 = 14'b10001000110111;
9'd229   : cube_lut_2 = 14'b10001000111010;
9'd230   : cube_lut_2 = 14'b10001000111100;
9'd231   : cube_lut_2 = 14'b10001000111110;
9'd232   : cube_lut_2 = 14'b10001001000001;
9'd233   : cube_lut_2 = 14'b10001001000011;
9'd234   : cube_lut_2 = 14'b10001001000101;
9'd235   : cube_lut_2 = 14'b10001001001000;
9'd236   : cube_lut_2 = 14'b10001001001010;
9'd237   : cube_lut_2 = 14'b10001001001100;
9'd238   : cube_lut_2 = 14'b10001001001111;
9'd239   : cube_lut_2 = 14'b10001001010001;
9'd240   : cube_lut_2 = 14'b10001001010011;
9'd241   : cube_lut_2 = 14'b10001001010101;
9'd242   : cube_lut_2 = 14'b10001001011000;
9'd243   : cube_lut_2 = 14'b10001001011010;
9'd244   : cube_lut_2 = 14'b10001001011100;
9'd245   : cube_lut_2 = 14'b10001001011111;
9'd246   : cube_lut_2 = 14'b10001001100001;
9'd247   : cube_lut_2 = 14'b10001001100011;
9'd248   : cube_lut_2 = 14'b10001001100110;
9'd249   : cube_lut_2 = 14'b10001001101000;
9'd250   : cube_lut_2 = 14'b10001001101010;
9'd251   : cube_lut_2 = 14'b10001001101101;
9'd252   : cube_lut_2 = 14'b10001001101111;
9'd253   : cube_lut_2 = 14'b10001001110001;
9'd254   : cube_lut_2 = 14'b10001001110011;
9'd255   : cube_lut_2 = 14'b10001001110110;
9'd256   : cube_lut_2 = 14'b10001001111000;
9'd257   : cube_lut_2 = 14'b10001001111010;
9'd258   : cube_lut_2 = 14'b10001001111101;
9'd259   : cube_lut_2 = 14'b10001001111111;
9'd260   : cube_lut_2 = 14'b10001010000001;
9'd261   : cube_lut_2 = 14'b10001010000100;
9'd262   : cube_lut_2 = 14'b10001010000110;
9'd263   : cube_lut_2 = 14'b10001010001000;
9'd264   : cube_lut_2 = 14'b10001010001010;
9'd265   : cube_lut_2 = 14'b10001010001101;
9'd266   : cube_lut_2 = 14'b10001010001111;
9'd267   : cube_lut_2 = 14'b10001010010001;
9'd268   : cube_lut_2 = 14'b10001010010100;
9'd269   : cube_lut_2 = 14'b10001010010110;
9'd270   : cube_lut_2 = 14'b10001010011000;
9'd271   : cube_lut_2 = 14'b10001010011010;
9'd272   : cube_lut_2 = 14'b10001010011101;
9'd273   : cube_lut_2 = 14'b10001010011111;
9'd274   : cube_lut_2 = 14'b10001010100001;
9'd275   : cube_lut_2 = 14'b10001010100100;
9'd276   : cube_lut_2 = 14'b10001010100110;
9'd277   : cube_lut_2 = 14'b10001010101000;
9'd278   : cube_lut_2 = 14'b10001010101010;
9'd279   : cube_lut_2 = 14'b10001010101101;
9'd280   : cube_lut_2 = 14'b10001010101111;
9'd281   : cube_lut_2 = 14'b10001010110001;
9'd282   : cube_lut_2 = 14'b10001010110011;
9'd283   : cube_lut_2 = 14'b10001010110110;
9'd284   : cube_lut_2 = 14'b10001010111000;
9'd285   : cube_lut_2 = 14'b10001010111010;
9'd286   : cube_lut_2 = 14'b10001010111100;
9'd287   : cube_lut_2 = 14'b10001010111111;
9'd288   : cube_lut_2 = 14'b10001011000001;
9'd289   : cube_lut_2 = 14'b10001011000011;
9'd290   : cube_lut_2 = 14'b10001011000110;
9'd291   : cube_lut_2 = 14'b10001011001000;
9'd292   : cube_lut_2 = 14'b10001011001010;
9'd293   : cube_lut_2 = 14'b10001011001100;
9'd294   : cube_lut_2 = 14'b10001011001111;
9'd295   : cube_lut_2 = 14'b10001011010001;
9'd296   : cube_lut_2 = 14'b10001011010011;
9'd297   : cube_lut_2 = 14'b10001011010101;
9'd298   : cube_lut_2 = 14'b10001011011000;
9'd299   : cube_lut_2 = 14'b10001011011010;
9'd300   : cube_lut_2 = 14'b10001011011100;
9'd301   : cube_lut_2 = 14'b10001011011110;
9'd302   : cube_lut_2 = 14'b10001011100001;
9'd303   : cube_lut_2 = 14'b10001011100011;
9'd304   : cube_lut_2 = 14'b10001011100101;
9'd305   : cube_lut_2 = 14'b10001011100111;
9'd306   : cube_lut_2 = 14'b10001011101010;
9'd307   : cube_lut_2 = 14'b10001011101100;
9'd308   : cube_lut_2 = 14'b10001011101110;
9'd309   : cube_lut_2 = 14'b10001011110000;
9'd310   : cube_lut_2 = 14'b10001011110010;
9'd311   : cube_lut_2 = 14'b10001011110101;
9'd312   : cube_lut_2 = 14'b10001011110111;
9'd313   : cube_lut_2 = 14'b10001011111001;
9'd314   : cube_lut_2 = 14'b10001011111011;
9'd315   : cube_lut_2 = 14'b10001011111110;
9'd316   : cube_lut_2 = 14'b10001100000000;
9'd317   : cube_lut_2 = 14'b10001100000010;
9'd318   : cube_lut_2 = 14'b10001100000100;
9'd319   : cube_lut_2 = 14'b10001100000111;
9'd320   : cube_lut_2 = 14'b10001100001001;
9'd321   : cube_lut_2 = 14'b10001100001011;
9'd322   : cube_lut_2 = 14'b10001100001101;
9'd323   : cube_lut_2 = 14'b10001100001111;
9'd324   : cube_lut_2 = 14'b10001100010010;
9'd325   : cube_lut_2 = 14'b10001100010100;
9'd326   : cube_lut_2 = 14'b10001100010110;
9'd327   : cube_lut_2 = 14'b10001100011000;
9'd328   : cube_lut_2 = 14'b10001100011011;
9'd329   : cube_lut_2 = 14'b10001100011101;
9'd330   : cube_lut_2 = 14'b10001100011111;
9'd331   : cube_lut_2 = 14'b10001100100001;
9'd332   : cube_lut_2 = 14'b10001100100011;
9'd333   : cube_lut_2 = 14'b10001100100110;
9'd334   : cube_lut_2 = 14'b10001100101000;
9'd335   : cube_lut_2 = 14'b10001100101010;
9'd336   : cube_lut_2 = 14'b10001100101100;
9'd337   : cube_lut_2 = 14'b10001100101110;
9'd338   : cube_lut_2 = 14'b10001100110001;
9'd339   : cube_lut_2 = 14'b10001100110011;
9'd340   : cube_lut_2 = 14'b10001100110101;
9'd341   : cube_lut_2 = 14'b10001100110111;
9'd342   : cube_lut_2 = 14'b10001100111001;
9'd343   : cube_lut_2 = 14'b10001100111100;
9'd344   : cube_lut_2 = 14'b10001100111110;
9'd345   : cube_lut_2 = 14'b10001101000000;
9'd346   : cube_lut_2 = 14'b10001101000010;
9'd347   : cube_lut_2 = 14'b10001101000100;
9'd348   : cube_lut_2 = 14'b10001101000111;
9'd349   : cube_lut_2 = 14'b10001101001001;
9'd350   : cube_lut_2 = 14'b10001101001011;
9'd351   : cube_lut_2 = 14'b10001101001101;
9'd352   : cube_lut_2 = 14'b10001101001111;
9'd353   : cube_lut_2 = 14'b10001101010010;
9'd354   : cube_lut_2 = 14'b10001101010100;
9'd355   : cube_lut_2 = 14'b10001101010110;
9'd356   : cube_lut_2 = 14'b10001101011000;
9'd357   : cube_lut_2 = 14'b10001101011010;
9'd358   : cube_lut_2 = 14'b10001101011101;
9'd359   : cube_lut_2 = 14'b10001101011111;
9'd360   : cube_lut_2 = 14'b10001101100001;
9'd361   : cube_lut_2 = 14'b10001101100011;
9'd362   : cube_lut_2 = 14'b10001101100101;
9'd363   : cube_lut_2 = 14'b10001101100111;
9'd364   : cube_lut_2 = 14'b10001101101010;
9'd365   : cube_lut_2 = 14'b10001101101100;
9'd366   : cube_lut_2 = 14'b10001101101110;
9'd367   : cube_lut_2 = 14'b10001101110000;
9'd368   : cube_lut_2 = 14'b10001101110010;
9'd369   : cube_lut_2 = 14'b10001101110100;
9'd370   : cube_lut_2 = 14'b10001101110111;
9'd371   : cube_lut_2 = 14'b10001101111001;
9'd372   : cube_lut_2 = 14'b10001101111011;
9'd373   : cube_lut_2 = 14'b10001101111101;
9'd374   : cube_lut_2 = 14'b10001101111111;
9'd375   : cube_lut_2 = 14'b10001110000001;
9'd376   : cube_lut_2 = 14'b10001110000100;
9'd377   : cube_lut_2 = 14'b10001110000110;
9'd378   : cube_lut_2 = 14'b10001110001000;
9'd379   : cube_lut_2 = 14'b10001110001010;
9'd380   : cube_lut_2 = 14'b10001110001100;
9'd381   : cube_lut_2 = 14'b10001110001110;
9'd382   : cube_lut_2 = 14'b10001110010001;
9'd383   : cube_lut_2 = 14'b10001110010011;
9'd384   : cube_lut_2 = 14'b10001110010101;
9'd385   : cube_lut_2 = 14'b10001110010111;
9'd386   : cube_lut_2 = 14'b10001110011001;
9'd387   : cube_lut_2 = 14'b10001110011011;
9'd388   : cube_lut_2 = 14'b10001110011110;
9'd389   : cube_lut_2 = 14'b10001110100000;
9'd390   : cube_lut_2 = 14'b10001110100010;
9'd391   : cube_lut_2 = 14'b10001110100100;
9'd392   : cube_lut_2 = 14'b10001110100110;
9'd393   : cube_lut_2 = 14'b10001110101000;
9'd394   : cube_lut_2 = 14'b10001110101010;
9'd395   : cube_lut_2 = 14'b10001110101101;
9'd396   : cube_lut_2 = 14'b10001110101111;
9'd397   : cube_lut_2 = 14'b10001110110001;
9'd398   : cube_lut_2 = 14'b10001110110011;
9'd399   : cube_lut_2 = 14'b10001110110101;
9'd400   : cube_lut_2 = 14'b10001110110111;
9'd401   : cube_lut_2 = 14'b10001110111001;
9'd402   : cube_lut_2 = 14'b10001110111100;
9'd403   : cube_lut_2 = 14'b10001110111110;
9'd404   : cube_lut_2 = 14'b10001111000000;
9'd405   : cube_lut_2 = 14'b10001111000010;
9'd406   : cube_lut_2 = 14'b10001111000100;
9'd407   : cube_lut_2 = 14'b10001111000110;
9'd408   : cube_lut_2 = 14'b10001111001000;
9'd409   : cube_lut_2 = 14'b10001111001011;
9'd410   : cube_lut_2 = 14'b10001111001101;
9'd411   : cube_lut_2 = 14'b10001111001111;
9'd412   : cube_lut_2 = 14'b10001111010001;
9'd413   : cube_lut_2 = 14'b10001111010011;
9'd414   : cube_lut_2 = 14'b10001111010101;
9'd415   : cube_lut_2 = 14'b10001111010111;
9'd416   : cube_lut_2 = 14'b10001111011001;
9'd417   : cube_lut_2 = 14'b10001111011100;
9'd418   : cube_lut_2 = 14'b10001111011110;
9'd419   : cube_lut_2 = 14'b10001111100000;
9'd420   : cube_lut_2 = 14'b10001111100010;
9'd421   : cube_lut_2 = 14'b10001111100100;
9'd422   : cube_lut_2 = 14'b10001111100110;
9'd423   : cube_lut_2 = 14'b10001111101000;
9'd424   : cube_lut_2 = 14'b10001111101010;
9'd425   : cube_lut_2 = 14'b10001111101100;
9'd426   : cube_lut_2 = 14'b10001111101111;
9'd427   : cube_lut_2 = 14'b10001111110001;
9'd428   : cube_lut_2 = 14'b10001111110011;
9'd429   : cube_lut_2 = 14'b10001111110101;
9'd430   : cube_lut_2 = 14'b10001111110111;
9'd431   : cube_lut_2 = 14'b10001111111001;
9'd432   : cube_lut_2 = 14'b10001111111011;
9'd433   : cube_lut_2 = 14'b10001111111101;
9'd434   : cube_lut_2 = 14'b10010000000000;
9'd435   : cube_lut_2 = 14'b10010000000010;
9'd436   : cube_lut_2 = 14'b10010000000100;
9'd437   : cube_lut_2 = 14'b10010000000110;
9'd438   : cube_lut_2 = 14'b10010000001000;
9'd439   : cube_lut_2 = 14'b10010000001010;
9'd440   : cube_lut_2 = 14'b10010000001100;
9'd441   : cube_lut_2 = 14'b10010000001110;
9'd442   : cube_lut_2 = 14'b10010000010000;
9'd443   : cube_lut_2 = 14'b10010000010010;
9'd444   : cube_lut_2 = 14'b10010000010101;
9'd445   : cube_lut_2 = 14'b10010000010111;
9'd446   : cube_lut_2 = 14'b10010000011001;
9'd447   : cube_lut_2 = 14'b10010000011011;
9'd448   : cube_lut_2 = 14'b10010000011101;
9'd449   : cube_lut_2 = 14'b10010000011111;
9'd450   : cube_lut_2 = 14'b10010000100001;
9'd451   : cube_lut_2 = 14'b10010000100011;
9'd452   : cube_lut_2 = 14'b10010000100101;
9'd453   : cube_lut_2 = 14'b10010000100111;
9'd454   : cube_lut_2 = 14'b10010000101001;
9'd455   : cube_lut_2 = 14'b10010000101100;
9'd456   : cube_lut_2 = 14'b10010000101110;
9'd457   : cube_lut_2 = 14'b10010000110000;
9'd458   : cube_lut_2 = 14'b10010000110010;
9'd459   : cube_lut_2 = 14'b10010000110100;
9'd460   : cube_lut_2 = 14'b10010000110110;
9'd461   : cube_lut_2 = 14'b10010000111000;
9'd462   : cube_lut_2 = 14'b10010000111010;
9'd463   : cube_lut_2 = 14'b10010000111100;
9'd464   : cube_lut_2 = 14'b10010000111110;
9'd465   : cube_lut_2 = 14'b10010001000000;
9'd466   : cube_lut_2 = 14'b10010001000010;
9'd467   : cube_lut_2 = 14'b10010001000101;
9'd468   : cube_lut_2 = 14'b10010001000111;
9'd469   : cube_lut_2 = 14'b10010001001001;
9'd470   : cube_lut_2 = 14'b10010001001011;
9'd471   : cube_lut_2 = 14'b10010001001101;
9'd472   : cube_lut_2 = 14'b10010001001111;
9'd473   : cube_lut_2 = 14'b10010001010001;
9'd474   : cube_lut_2 = 14'b10010001010011;
9'd475   : cube_lut_2 = 14'b10010001010101;
9'd476   : cube_lut_2 = 14'b10010001010111;
9'd477   : cube_lut_2 = 14'b10010001011001;
9'd478   : cube_lut_2 = 14'b10010001011011;
9'd479   : cube_lut_2 = 14'b10010001011101;
9'd480   : cube_lut_2 = 14'b10010001011111;
9'd481   : cube_lut_2 = 14'b10010001100001;
9'd482   : cube_lut_2 = 14'b10010001100100;
9'd483   : cube_lut_2 = 14'b10010001100110;
9'd484   : cube_lut_2 = 14'b10010001101000;
9'd485   : cube_lut_2 = 14'b10010001101010;
9'd486   : cube_lut_2 = 14'b10010001101100;
9'd487   : cube_lut_2 = 14'b10010001101110;
9'd488   : cube_lut_2 = 14'b10010001110000;
9'd489   : cube_lut_2 = 14'b10010001110010;
9'd490   : cube_lut_2 = 14'b10010001110100;
9'd491   : cube_lut_2 = 14'b10010001110110;
9'd492   : cube_lut_2 = 14'b10010001111000;
9'd493   : cube_lut_2 = 14'b10010001111010;
9'd494   : cube_lut_2 = 14'b10010001111100;
9'd495   : cube_lut_2 = 14'b10010001111110;
9'd496   : cube_lut_2 = 14'b10010010000000;
9'd497   : cube_lut_2 = 14'b10010010000010;
9'd498   : cube_lut_2 = 14'b10010010000100;
9'd499   : cube_lut_2 = 14'b10010010000110;
9'd500   : cube_lut_2 = 14'b10010010001001;
9'd501   : cube_lut_2 = 14'b10010010001011;
9'd502   : cube_lut_2 = 14'b10010010001101;
9'd503   : cube_lut_2 = 14'b10010010001111;
9'd504   : cube_lut_2 = 14'b10010010010001;
9'd505   : cube_lut_2 = 14'b10010010010011;
9'd506   : cube_lut_2 = 14'b10010010010101;
9'd507   : cube_lut_2 = 14'b10010010010111;
9'd508   : cube_lut_2 = 14'b10010010011001;
9'd509   : cube_lut_2 = 14'b10010010011011;
9'd510   : cube_lut_2 = 14'b10010010011101;
9'd511   : cube_lut_2 = 14'b10010010011111;

    endcase
end

always@* begin
    
    cube_lut_3 = 0;
    
    case(i_data[8:0])
 
 9'd0   : cube_lut_3 = 14'b10010010100001;
9'd1   : cube_lut_3 = 14'b10010010100011;
9'd2   : cube_lut_3 = 14'b10010010100101;
9'd3   : cube_lut_3 = 14'b10010010100111;
9'd4   : cube_lut_3 = 14'b10010010101001;
9'd5   : cube_lut_3 = 14'b10010010101011;
9'd6   : cube_lut_3 = 14'b10010010101101;
9'd7   : cube_lut_3 = 14'b10010010101111;
9'd8   : cube_lut_3 = 14'b10010010110001;
9'd9   : cube_lut_3 = 14'b10010010110011;
9'd10   : cube_lut_3 = 14'b10010010110101;
9'd11   : cube_lut_3 = 14'b10010010110111;
9'd12   : cube_lut_3 = 14'b10010010111001;
9'd13   : cube_lut_3 = 14'b10010010111011;
9'd14   : cube_lut_3 = 14'b10010010111101;
9'd15   : cube_lut_3 = 14'b10010010111111;
9'd16   : cube_lut_3 = 14'b10010011000001;
9'd17   : cube_lut_3 = 14'b10010011000011;
9'd18   : cube_lut_3 = 14'b10010011000101;
9'd19   : cube_lut_3 = 14'b10010011001000;
9'd20   : cube_lut_3 = 14'b10010011001010;
9'd21   : cube_lut_3 = 14'b10010011001100;
9'd22   : cube_lut_3 = 14'b10010011001110;
9'd23   : cube_lut_3 = 14'b10010011010000;
9'd24   : cube_lut_3 = 14'b10010011010010;
9'd25   : cube_lut_3 = 14'b10010011010100;
9'd26   : cube_lut_3 = 14'b10010011010110;
9'd27   : cube_lut_3 = 14'b10010011011000;
9'd28   : cube_lut_3 = 14'b10010011011010;
9'd29   : cube_lut_3 = 14'b10010011011100;
9'd30   : cube_lut_3 = 14'b10010011011110;
9'd31   : cube_lut_3 = 14'b10010011100000;
9'd32   : cube_lut_3 = 14'b10010011100010;
9'd33   : cube_lut_3 = 14'b10010011100100;
9'd34   : cube_lut_3 = 14'b10010011100110;
9'd35   : cube_lut_3 = 14'b10010011101000;
9'd36   : cube_lut_3 = 14'b10010011101010;
9'd37   : cube_lut_3 = 14'b10010011101100;
9'd38   : cube_lut_3 = 14'b10010011101110;
9'd39   : cube_lut_3 = 14'b10010011110000;
9'd40   : cube_lut_3 = 14'b10010011110010;
9'd41   : cube_lut_3 = 14'b10010011110100;
9'd42   : cube_lut_3 = 14'b10010011110110;
9'd43   : cube_lut_3 = 14'b10010011111000;
9'd44   : cube_lut_3 = 14'b10010011111010;
9'd45   : cube_lut_3 = 14'b10010011111100;
9'd46   : cube_lut_3 = 14'b10010011111110;
9'd47   : cube_lut_3 = 14'b10010100000000;
9'd48   : cube_lut_3 = 14'b10010100000010;
9'd49   : cube_lut_3 = 14'b10010100000100;
9'd50   : cube_lut_3 = 14'b10010100000110;
9'd51   : cube_lut_3 = 14'b10010100001000;
9'd52   : cube_lut_3 = 14'b10010100001010;
9'd53   : cube_lut_3 = 14'b10010100001100;
9'd54   : cube_lut_3 = 14'b10010100001110;
9'd55   : cube_lut_3 = 14'b10010100010000;
9'd56   : cube_lut_3 = 14'b10010100010010;
9'd57   : cube_lut_3 = 14'b10010100010100;
9'd58   : cube_lut_3 = 14'b10010100010110;
9'd59   : cube_lut_3 = 14'b10010100011000;
9'd60   : cube_lut_3 = 14'b10010100011010;
9'd61   : cube_lut_3 = 14'b10010100011100;
9'd62   : cube_lut_3 = 14'b10010100011110;
9'd63   : cube_lut_3 = 14'b10010100011111;
9'd64   : cube_lut_3 = 14'b10010100100001;
9'd65   : cube_lut_3 = 14'b10010100100011;
9'd66   : cube_lut_3 = 14'b10010100100101;
9'd67   : cube_lut_3 = 14'b10010100100111;
9'd68   : cube_lut_3 = 14'b10010100101001;
9'd69   : cube_lut_3 = 14'b10010100101011;
9'd70   : cube_lut_3 = 14'b10010100101101;
9'd71   : cube_lut_3 = 14'b10010100101111;
9'd72   : cube_lut_3 = 14'b10010100110001;
9'd73   : cube_lut_3 = 14'b10010100110011;
9'd74   : cube_lut_3 = 14'b10010100110101;
9'd75   : cube_lut_3 = 14'b10010100110111;
9'd76   : cube_lut_3 = 14'b10010100111001;
9'd77   : cube_lut_3 = 14'b10010100111011;
9'd78   : cube_lut_3 = 14'b10010100111101;
9'd79   : cube_lut_3 = 14'b10010100111111;
9'd80   : cube_lut_3 = 14'b10010101000001;
9'd81   : cube_lut_3 = 14'b10010101000011;
9'd82   : cube_lut_3 = 14'b10010101000101;
9'd83   : cube_lut_3 = 14'b10010101000111;
9'd84   : cube_lut_3 = 14'b10010101001001;
9'd85   : cube_lut_3 = 14'b10010101001011;
9'd86   : cube_lut_3 = 14'b10010101001101;
9'd87   : cube_lut_3 = 14'b10010101001111;
9'd88   : cube_lut_3 = 14'b10010101010001;
9'd89   : cube_lut_3 = 14'b10010101010011;
9'd90   : cube_lut_3 = 14'b10010101010101;
9'd91   : cube_lut_3 = 14'b10010101010111;
9'd92   : cube_lut_3 = 14'b10010101011001;
9'd93   : cube_lut_3 = 14'b10010101011011;
9'd94   : cube_lut_3 = 14'b10010101011101;
9'd95   : cube_lut_3 = 14'b10010101011110;
9'd96   : cube_lut_3 = 14'b10010101100000;
9'd97   : cube_lut_3 = 14'b10010101100010;
9'd98   : cube_lut_3 = 14'b10010101100100;
9'd99   : cube_lut_3 = 14'b10010101100110;
9'd100   : cube_lut_3 = 14'b10010101101000;
9'd101   : cube_lut_3 = 14'b10010101101010;
9'd102   : cube_lut_3 = 14'b10010101101100;
9'd103   : cube_lut_3 = 14'b10010101101110;
9'd104   : cube_lut_3 = 14'b10010101110000;
9'd105   : cube_lut_3 = 14'b10010101110010;
9'd106   : cube_lut_3 = 14'b10010101110100;
9'd107   : cube_lut_3 = 14'b10010101110110;
9'd108   : cube_lut_3 = 14'b10010101111000;
9'd109   : cube_lut_3 = 14'b10010101111010;
9'd110   : cube_lut_3 = 14'b10010101111100;
9'd111   : cube_lut_3 = 14'b10010101111110;
9'd112   : cube_lut_3 = 14'b10010110000000;
9'd113   : cube_lut_3 = 14'b10010110000010;
9'd114   : cube_lut_3 = 14'b10010110000011;
9'd115   : cube_lut_3 = 14'b10010110000101;
9'd116   : cube_lut_3 = 14'b10010110000111;
9'd117   : cube_lut_3 = 14'b10010110001001;
9'd118   : cube_lut_3 = 14'b10010110001011;
9'd119   : cube_lut_3 = 14'b10010110001101;
9'd120   : cube_lut_3 = 14'b10010110001111;
9'd121   : cube_lut_3 = 14'b10010110010001;
9'd122   : cube_lut_3 = 14'b10010110010011;
9'd123   : cube_lut_3 = 14'b10010110010101;
9'd124   : cube_lut_3 = 14'b10010110010111;
9'd125   : cube_lut_3 = 14'b10010110011001;
9'd126   : cube_lut_3 = 14'b10010110011011;
9'd127   : cube_lut_3 = 14'b10010110011101;
9'd128   : cube_lut_3 = 14'b10010110011111;
9'd129   : cube_lut_3 = 14'b10010110100000;
9'd130   : cube_lut_3 = 14'b10010110100010;
9'd131   : cube_lut_3 = 14'b10010110100100;
9'd132   : cube_lut_3 = 14'b10010110100110;
9'd133   : cube_lut_3 = 14'b10010110101000;
9'd134   : cube_lut_3 = 14'b10010110101010;
9'd135   : cube_lut_3 = 14'b10010110101100;
9'd136   : cube_lut_3 = 14'b10010110101110;
9'd137   : cube_lut_3 = 14'b10010110110000;
9'd138   : cube_lut_3 = 14'b10010110110010;
9'd139   : cube_lut_3 = 14'b10010110110100;
9'd140   : cube_lut_3 = 14'b10010110110110;
9'd141   : cube_lut_3 = 14'b10010110111000;
9'd142   : cube_lut_3 = 14'b10010110111010;
9'd143   : cube_lut_3 = 14'b10010110111011;
9'd144   : cube_lut_3 = 14'b10010110111101;
9'd145   : cube_lut_3 = 14'b10010110111111;
9'd146   : cube_lut_3 = 14'b10010111000001;
9'd147   : cube_lut_3 = 14'b10010111000011;
9'd148   : cube_lut_3 = 14'b10010111000101;
9'd149   : cube_lut_3 = 14'b10010111000111;
9'd150   : cube_lut_3 = 14'b10010111001001;
9'd151   : cube_lut_3 = 14'b10010111001011;
9'd152   : cube_lut_3 = 14'b10010111001101;
9'd153   : cube_lut_3 = 14'b10010111001111;
9'd154   : cube_lut_3 = 14'b10010111010000;
9'd155   : cube_lut_3 = 14'b10010111010010;
9'd156   : cube_lut_3 = 14'b10010111010100;
9'd157   : cube_lut_3 = 14'b10010111010110;
9'd158   : cube_lut_3 = 14'b10010111011000;
9'd159   : cube_lut_3 = 14'b10010111011010;
9'd160   : cube_lut_3 = 14'b10010111011100;
9'd161   : cube_lut_3 = 14'b10010111011110;
9'd162   : cube_lut_3 = 14'b10010111100000;
9'd163   : cube_lut_3 = 14'b10010111100010;
9'd164   : cube_lut_3 = 14'b10010111100100;
9'd165   : cube_lut_3 = 14'b10010111100101;
9'd166   : cube_lut_3 = 14'b10010111100111;
9'd167   : cube_lut_3 = 14'b10010111101001;
9'd168   : cube_lut_3 = 14'b10010111101011;
9'd169   : cube_lut_3 = 14'b10010111101101;
9'd170   : cube_lut_3 = 14'b10010111101111;
9'd171   : cube_lut_3 = 14'b10010111110001;
9'd172   : cube_lut_3 = 14'b10010111110011;
9'd173   : cube_lut_3 = 14'b10010111110101;
9'd174   : cube_lut_3 = 14'b10010111110111;
9'd175   : cube_lut_3 = 14'b10010111111000;
9'd176   : cube_lut_3 = 14'b10010111111010;
9'd177   : cube_lut_3 = 14'b10010111111100;
9'd178   : cube_lut_3 = 14'b10010111111110;
9'd179   : cube_lut_3 = 14'b10011000000000;
9'd180   : cube_lut_3 = 14'b10011000000010;
9'd181   : cube_lut_3 = 14'b10011000000100;
9'd182   : cube_lut_3 = 14'b10011000000110;
9'd183   : cube_lut_3 = 14'b10011000001000;
9'd184   : cube_lut_3 = 14'b10011000001001;
9'd185   : cube_lut_3 = 14'b10011000001011;
9'd186   : cube_lut_3 = 14'b10011000001101;
9'd187   : cube_lut_3 = 14'b10011000001111;
9'd188   : cube_lut_3 = 14'b10011000010001;
9'd189   : cube_lut_3 = 14'b10011000010011;
9'd190   : cube_lut_3 = 14'b10011000010101;
9'd191   : cube_lut_3 = 14'b10011000010111;
9'd192   : cube_lut_3 = 14'b10011000011000;
9'd193   : cube_lut_3 = 14'b10011000011010;
9'd194   : cube_lut_3 = 14'b10011000011100;
9'd195   : cube_lut_3 = 14'b10011000011110;
9'd196   : cube_lut_3 = 14'b10011000100000;
9'd197   : cube_lut_3 = 14'b10011000100010;
9'd198   : cube_lut_3 = 14'b10011000100100;
9'd199   : cube_lut_3 = 14'b10011000100110;
9'd200   : cube_lut_3 = 14'b10011000101000;
9'd201   : cube_lut_3 = 14'b10011000101001;
9'd202   : cube_lut_3 = 14'b10011000101011;
9'd203   : cube_lut_3 = 14'b10011000101101;
9'd204   : cube_lut_3 = 14'b10011000101111;
9'd205   : cube_lut_3 = 14'b10011000110001;
9'd206   : cube_lut_3 = 14'b10011000110011;
9'd207   : cube_lut_3 = 14'b10011000110101;
9'd208   : cube_lut_3 = 14'b10011000110111;
9'd209   : cube_lut_3 = 14'b10011000111000;
9'd210   : cube_lut_3 = 14'b10011000111010;
9'd211   : cube_lut_3 = 14'b10011000111100;
9'd212   : cube_lut_3 = 14'b10011000111110;
9'd213   : cube_lut_3 = 14'b10011001000000;
9'd214   : cube_lut_3 = 14'b10011001000010;
9'd215   : cube_lut_3 = 14'b10011001000100;
9'd216   : cube_lut_3 = 14'b10011001000101;
9'd217   : cube_lut_3 = 14'b10011001000111;
9'd218   : cube_lut_3 = 14'b10011001001001;
9'd219   : cube_lut_3 = 14'b10011001001011;
9'd220   : cube_lut_3 = 14'b10011001001101;
9'd221   : cube_lut_3 = 14'b10011001001111;
9'd222   : cube_lut_3 = 14'b10011001010001;
9'd223   : cube_lut_3 = 14'b10011001010010;
9'd224   : cube_lut_3 = 14'b10011001010100;
9'd225   : cube_lut_3 = 14'b10011001010110;
9'd226   : cube_lut_3 = 14'b10011001011000;
9'd227   : cube_lut_3 = 14'b10011001011010;
9'd228   : cube_lut_3 = 14'b10011001011100;
9'd229   : cube_lut_3 = 14'b10011001011110;
9'd230   : cube_lut_3 = 14'b10011001011111;
9'd231   : cube_lut_3 = 14'b10011001100001;
9'd232   : cube_lut_3 = 14'b10011001100011;
9'd233   : cube_lut_3 = 14'b10011001100101;
9'd234   : cube_lut_3 = 14'b10011001100111;
9'd235   : cube_lut_3 = 14'b10011001101001;
9'd236   : cube_lut_3 = 14'b10011001101011;
9'd237   : cube_lut_3 = 14'b10011001101100;
9'd238   : cube_lut_3 = 14'b10011001101110;
9'd239   : cube_lut_3 = 14'b10011001110000;
9'd240   : cube_lut_3 = 14'b10011001110010;
9'd241   : cube_lut_3 = 14'b10011001110100;
9'd242   : cube_lut_3 = 14'b10011001110110;
9'd243   : cube_lut_3 = 14'b10011001111000;
9'd244   : cube_lut_3 = 14'b10011001111001;
9'd245   : cube_lut_3 = 14'b10011001111011;
9'd246   : cube_lut_3 = 14'b10011001111101;
9'd247   : cube_lut_3 = 14'b10011001111111;
9'd248   : cube_lut_3 = 14'b10011010000001;
9'd249   : cube_lut_3 = 14'b10011010000011;
9'd250   : cube_lut_3 = 14'b10011010000100;
9'd251   : cube_lut_3 = 14'b10011010000110;
9'd252   : cube_lut_3 = 14'b10011010001000;
9'd253   : cube_lut_3 = 14'b10011010001010;
9'd254   : cube_lut_3 = 14'b10011010001100;
9'd255   : cube_lut_3 = 14'b10011010001110;
9'd256   : cube_lut_3 = 14'b10011010001111;
9'd257   : cube_lut_3 = 14'b10011010010001;
9'd258   : cube_lut_3 = 14'b10011010010011;
9'd259   : cube_lut_3 = 14'b10011010010101;
9'd260   : cube_lut_3 = 14'b10011010010111;
9'd261   : cube_lut_3 = 14'b10011010011001;
9'd262   : cube_lut_3 = 14'b10011010011010;
9'd263   : cube_lut_3 = 14'b10011010011100;
9'd264   : cube_lut_3 = 14'b10011010011110;
9'd265   : cube_lut_3 = 14'b10011010100000;
9'd266   : cube_lut_3 = 14'b10011010100010;
9'd267   : cube_lut_3 = 14'b10011010100100;
9'd268   : cube_lut_3 = 14'b10011010100101;
9'd269   : cube_lut_3 = 14'b10011010100111;
9'd270   : cube_lut_3 = 14'b10011010101001;
9'd271   : cube_lut_3 = 14'b10011010101011;
9'd272   : cube_lut_3 = 14'b10011010101101;
9'd273   : cube_lut_3 = 14'b10011010101111;
9'd274   : cube_lut_3 = 14'b10011010110000;
9'd275   : cube_lut_3 = 14'b10011010110010;
9'd276   : cube_lut_3 = 14'b10011010110100;
9'd277   : cube_lut_3 = 14'b10011010110110;
9'd278   : cube_lut_3 = 14'b10011010111000;
9'd279   : cube_lut_3 = 14'b10011010111001;
9'd280   : cube_lut_3 = 14'b10011010111011;
9'd281   : cube_lut_3 = 14'b10011010111101;
9'd282   : cube_lut_3 = 14'b10011010111111;
9'd283   : cube_lut_3 = 14'b10011011000001;
9'd284   : cube_lut_3 = 14'b10011011000011;
9'd285   : cube_lut_3 = 14'b10011011000100;
9'd286   : cube_lut_3 = 14'b10011011000110;
9'd287   : cube_lut_3 = 14'b10011011001000;
9'd288   : cube_lut_3 = 14'b10011011001010;
9'd289   : cube_lut_3 = 14'b10011011001100;
9'd290   : cube_lut_3 = 14'b10011011001101;
9'd291   : cube_lut_3 = 14'b10011011001111;
9'd292   : cube_lut_3 = 14'b10011011010001;
9'd293   : cube_lut_3 = 14'b10011011010011;
9'd294   : cube_lut_3 = 14'b10011011010101;
9'd295   : cube_lut_3 = 14'b10011011010111;
9'd296   : cube_lut_3 = 14'b10011011011000;
9'd297   : cube_lut_3 = 14'b10011011011010;
9'd298   : cube_lut_3 = 14'b10011011011100;
9'd299   : cube_lut_3 = 14'b10011011011110;
9'd300   : cube_lut_3 = 14'b10011011100000;
9'd301   : cube_lut_3 = 14'b10011011100001;
9'd302   : cube_lut_3 = 14'b10011011100011;
9'd303   : cube_lut_3 = 14'b10011011100101;
9'd304   : cube_lut_3 = 14'b10011011100111;
9'd305   : cube_lut_3 = 14'b10011011101001;
9'd306   : cube_lut_3 = 14'b10011011101010;
9'd307   : cube_lut_3 = 14'b10011011101100;
9'd308   : cube_lut_3 = 14'b10011011101110;
9'd309   : cube_lut_3 = 14'b10011011110000;
9'd310   : cube_lut_3 = 14'b10011011110010;
9'd311   : cube_lut_3 = 14'b10011011110011;
9'd312   : cube_lut_3 = 14'b10011011110101;
9'd313   : cube_lut_3 = 14'b10011011110111;
9'd314   : cube_lut_3 = 14'b10011011111001;
9'd315   : cube_lut_3 = 14'b10011011111011;
9'd316   : cube_lut_3 = 14'b10011011111100;
9'd317   : cube_lut_3 = 14'b10011011111110;
9'd318   : cube_lut_3 = 14'b10011100000000;
9'd319   : cube_lut_3 = 14'b10011100000010;
9'd320   : cube_lut_3 = 14'b10011100000100;
9'd321   : cube_lut_3 = 14'b10011100000101;
9'd322   : cube_lut_3 = 14'b10011100000111;
9'd323   : cube_lut_3 = 14'b10011100001001;
9'd324   : cube_lut_3 = 14'b10011100001011;
9'd325   : cube_lut_3 = 14'b10011100001101;
9'd326   : cube_lut_3 = 14'b10011100001110;
9'd327   : cube_lut_3 = 14'b10011100010000;
9'd328   : cube_lut_3 = 14'b10011100010010;
9'd329   : cube_lut_3 = 14'b10011100010100;
9'd330   : cube_lut_3 = 14'b10011100010110;
9'd331   : cube_lut_3 = 14'b10011100010111;
9'd332   : cube_lut_3 = 14'b10011100011001;
9'd333   : cube_lut_3 = 14'b10011100011011;
9'd334   : cube_lut_3 = 14'b10011100011101;
9'd335   : cube_lut_3 = 14'b10011100011110;
9'd336   : cube_lut_3 = 14'b10011100100000;
9'd337   : cube_lut_3 = 14'b10011100100010;
9'd338   : cube_lut_3 = 14'b10011100100100;
9'd339   : cube_lut_3 = 14'b10011100100110;
9'd340   : cube_lut_3 = 14'b10011100100111;
9'd341   : cube_lut_3 = 14'b10011100101001;
9'd342   : cube_lut_3 = 14'b10011100101011;
9'd343   : cube_lut_3 = 14'b10011100101101;
9'd344   : cube_lut_3 = 14'b10011100101110;
9'd345   : cube_lut_3 = 14'b10011100110000;
9'd346   : cube_lut_3 = 14'b10011100110010;
9'd347   : cube_lut_3 = 14'b10011100110100;
9'd348   : cube_lut_3 = 14'b10011100110110;
9'd349   : cube_lut_3 = 14'b10011100110111;
9'd350   : cube_lut_3 = 14'b10011100111001;
9'd351   : cube_lut_3 = 14'b10011100111011;
9'd352   : cube_lut_3 = 14'b10011100111101;
9'd353   : cube_lut_3 = 14'b10011100111110;
9'd354   : cube_lut_3 = 14'b10011101000000;
9'd355   : cube_lut_3 = 14'b10011101000010;
9'd356   : cube_lut_3 = 14'b10011101000100;
9'd357   : cube_lut_3 = 14'b10011101000110;
9'd358   : cube_lut_3 = 14'b10011101000111;
9'd359   : cube_lut_3 = 14'b10011101001001;
9'd360   : cube_lut_3 = 14'b10011101001011;
9'd361   : cube_lut_3 = 14'b10011101001101;
9'd362   : cube_lut_3 = 14'b10011101001110;
9'd363   : cube_lut_3 = 14'b10011101010000;
9'd364   : cube_lut_3 = 14'b10011101010010;
9'd365   : cube_lut_3 = 14'b10011101010100;
9'd366   : cube_lut_3 = 14'b10011101010101;
9'd367   : cube_lut_3 = 14'b10011101010111;
9'd368   : cube_lut_3 = 14'b10011101011001;
9'd369   : cube_lut_3 = 14'b10011101011011;
9'd370   : cube_lut_3 = 14'b10011101011100;
9'd371   : cube_lut_3 = 14'b10011101011110;
9'd372   : cube_lut_3 = 14'b10011101100000;
9'd373   : cube_lut_3 = 14'b10011101100010;
9'd374   : cube_lut_3 = 14'b10011101100100;
9'd375   : cube_lut_3 = 14'b10011101100101;
9'd376   : cube_lut_3 = 14'b10011101100111;
9'd377   : cube_lut_3 = 14'b10011101101001;
9'd378   : cube_lut_3 = 14'b10011101101011;
9'd379   : cube_lut_3 = 14'b10011101101100;
9'd380   : cube_lut_3 = 14'b10011101101110;
9'd381   : cube_lut_3 = 14'b10011101110000;
9'd382   : cube_lut_3 = 14'b10011101110010;
9'd383   : cube_lut_3 = 14'b10011101110011;
9'd384   : cube_lut_3 = 14'b10011101110101;
9'd385   : cube_lut_3 = 14'b10011101110111;
9'd386   : cube_lut_3 = 14'b10011101111001;
9'd387   : cube_lut_3 = 14'b10011101111010;
9'd388   : cube_lut_3 = 14'b10011101111100;
9'd389   : cube_lut_3 = 14'b10011101111110;
9'd390   : cube_lut_3 = 14'b10011110000000;
9'd391   : cube_lut_3 = 14'b10011110000001;
9'd392   : cube_lut_3 = 14'b10011110000011;
9'd393   : cube_lut_3 = 14'b10011110000101;
9'd394   : cube_lut_3 = 14'b10011110000111;
9'd395   : cube_lut_3 = 14'b10011110001000;
9'd396   : cube_lut_3 = 14'b10011110001010;
9'd397   : cube_lut_3 = 14'b10011110001100;
9'd398   : cube_lut_3 = 14'b10011110001110;
9'd399   : cube_lut_3 = 14'b10011110001111;
9'd400   : cube_lut_3 = 14'b10011110010001;
9'd401   : cube_lut_3 = 14'b10011110010011;
9'd402   : cube_lut_3 = 14'b10011110010101;
9'd403   : cube_lut_3 = 14'b10011110010110;
9'd404   : cube_lut_3 = 14'b10011110011000;
9'd405   : cube_lut_3 = 14'b10011110011010;
9'd406   : cube_lut_3 = 14'b10011110011100;
9'd407   : cube_lut_3 = 14'b10011110011101;
9'd408   : cube_lut_3 = 14'b10011110011111;
9'd409   : cube_lut_3 = 14'b10011110100001;
9'd410   : cube_lut_3 = 14'b10011110100010;
9'd411   : cube_lut_3 = 14'b10011110100100;
9'd412   : cube_lut_3 = 14'b10011110100110;
9'd413   : cube_lut_3 = 14'b10011110101000;
9'd414   : cube_lut_3 = 14'b10011110101001;
9'd415   : cube_lut_3 = 14'b10011110101011;
9'd416   : cube_lut_3 = 14'b10011110101101;
9'd417   : cube_lut_3 = 14'b10011110101111;
9'd418   : cube_lut_3 = 14'b10011110110000;
9'd419   : cube_lut_3 = 14'b10011110110010;
9'd420   : cube_lut_3 = 14'b10011110110100;
9'd421   : cube_lut_3 = 14'b10011110110110;
9'd422   : cube_lut_3 = 14'b10011110110111;
9'd423   : cube_lut_3 = 14'b10011110111001;
9'd424   : cube_lut_3 = 14'b10011110111011;
9'd425   : cube_lut_3 = 14'b10011110111101;
9'd426   : cube_lut_3 = 14'b10011110111110;
9'd427   : cube_lut_3 = 14'b10011111000000;
9'd428   : cube_lut_3 = 14'b10011111000010;
9'd429   : cube_lut_3 = 14'b10011111000011;
9'd430   : cube_lut_3 = 14'b10011111000101;
9'd431   : cube_lut_3 = 14'b10011111000111;
9'd432   : cube_lut_3 = 14'b10011111001001;
9'd433   : cube_lut_3 = 14'b10011111001010;
9'd434   : cube_lut_3 = 14'b10011111001100;
9'd435   : cube_lut_3 = 14'b10011111001110;
9'd436   : cube_lut_3 = 14'b10011111001111;
9'd437   : cube_lut_3 = 14'b10011111010001;
9'd438   : cube_lut_3 = 14'b10011111010011;
9'd439   : cube_lut_3 = 14'b10011111010101;
9'd440   : cube_lut_3 = 14'b10011111010110;
9'd441   : cube_lut_3 = 14'b10011111011000;
9'd442   : cube_lut_3 = 14'b10011111011010;
9'd443   : cube_lut_3 = 14'b10011111011100;
9'd444   : cube_lut_3 = 14'b10011111011101;
9'd445   : cube_lut_3 = 14'b10011111011111;
9'd446   : cube_lut_3 = 14'b10011111100001;
9'd447   : cube_lut_3 = 14'b10011111100010;
9'd448   : cube_lut_3 = 14'b10011111100100;
9'd449   : cube_lut_3 = 14'b10011111100110;
9'd450   : cube_lut_3 = 14'b10011111101000;
9'd451   : cube_lut_3 = 14'b10011111101001;
9'd452   : cube_lut_3 = 14'b10011111101011;
9'd453   : cube_lut_3 = 14'b10011111101101;
9'd454   : cube_lut_3 = 14'b10011111101110;
9'd455   : cube_lut_3 = 14'b10011111110000;
9'd456   : cube_lut_3 = 14'b10011111110010;
9'd457   : cube_lut_3 = 14'b10011111110100;
9'd458   : cube_lut_3 = 14'b10011111110101;
9'd459   : cube_lut_3 = 14'b10011111110111;
9'd460   : cube_lut_3 = 14'b10011111111001;
9'd461   : cube_lut_3 = 14'b10011111111010;
9'd462   : cube_lut_3 = 14'b10011111111100;
9'd463   : cube_lut_3 = 14'b10011111111110;
9'd464   : cube_lut_3 = 14'b10100000000000;
9'd465   : cube_lut_3 = 14'b10100000000001;
9'd466   : cube_lut_3 = 14'b10100000000011;
9'd467   : cube_lut_3 = 14'b10100000000101;
9'd468   : cube_lut_3 = 14'b10100000000110;
9'd469   : cube_lut_3 = 14'b10100000001000;
9'd470   : cube_lut_3 = 14'b10100000001010;
9'd471   : cube_lut_3 = 14'b10100000001011;
9'd472   : cube_lut_3 = 14'b10100000001101;
9'd473   : cube_lut_3 = 14'b10100000001111;
9'd474   : cube_lut_3 = 14'b10100000010001;
9'd475   : cube_lut_3 = 14'b10100000010010;
9'd476   : cube_lut_3 = 14'b10100000010100;
9'd477   : cube_lut_3 = 14'b10100000010110;
9'd478   : cube_lut_3 = 14'b10100000010111;
9'd479   : cube_lut_3 = 14'b10100000011001;
9'd480   : cube_lut_3 = 14'b10100000011011;
9'd481   : cube_lut_3 = 14'b10100000011100;
9'd482   : cube_lut_3 = 14'b10100000011110;
9'd483   : cube_lut_3 = 14'b10100000100000;
9'd484   : cube_lut_3 = 14'b10100000100010;
9'd485   : cube_lut_3 = 14'b10100000100011;
9'd486   : cube_lut_3 = 14'b10100000100101;
9'd487   : cube_lut_3 = 14'b10100000100111;
9'd488   : cube_lut_3 = 14'b10100000101000;
9'd489   : cube_lut_3 = 14'b10100000101010;
9'd490   : cube_lut_3 = 14'b10100000101100;
9'd491   : cube_lut_3 = 14'b10100000101101;
9'd492   : cube_lut_3 = 14'b10100000101111;
9'd493   : cube_lut_3 = 14'b10100000110001;
9'd494   : cube_lut_3 = 14'b10100000110010;
9'd495   : cube_lut_3 = 14'b10100000110100;
9'd496   : cube_lut_3 = 14'b10100000110110;
9'd497   : cube_lut_3 = 14'b10100000111000;
9'd498   : cube_lut_3 = 14'b10100000111001;
9'd499   : cube_lut_3 = 14'b10100000111011;
9'd500   : cube_lut_3 = 14'b10100000111101;
9'd501   : cube_lut_3 = 14'b10100000111110;
9'd502   : cube_lut_3 = 14'b10100001000000;
9'd503   : cube_lut_3 = 14'b10100001000010;
9'd504   : cube_lut_3 = 14'b10100001000011;
9'd505   : cube_lut_3 = 14'b10100001000101;
9'd506   : cube_lut_3 = 14'b10100001000111;
9'd507   : cube_lut_3 = 14'b10100001001000;
9'd508   : cube_lut_3 = 14'b10100001001010;
9'd509   : cube_lut_3 = 14'b10100001001100;
9'd510   : cube_lut_3 = 14'b10100001001101;
9'd511   : cube_lut_3 = 14'b10100001001111;

    endcase
end

always@* begin
    
    cube_lut_4 = 0;
    
    case(i_data[8:0])
 
 9'd0   : cube_lut_4 = 14'b10100001010001;
9'd1   : cube_lut_4 = 14'b10100001010010;
9'd2   : cube_lut_4 = 14'b10100001010100;
9'd3   : cube_lut_4 = 14'b10100001010110;
9'd4   : cube_lut_4 = 14'b10100001010111;
9'd5   : cube_lut_4 = 14'b10100001011001;
9'd6   : cube_lut_4 = 14'b10100001011011;
9'd7   : cube_lut_4 = 14'b10100001011101;
9'd8   : cube_lut_4 = 14'b10100001011110;
9'd9   : cube_lut_4 = 14'b10100001100000;
9'd10   : cube_lut_4 = 14'b10100001100010;
9'd11   : cube_lut_4 = 14'b10100001100011;
9'd12   : cube_lut_4 = 14'b10100001100101;
9'd13   : cube_lut_4 = 14'b10100001100111;
9'd14   : cube_lut_4 = 14'b10100001101000;
9'd15   : cube_lut_4 = 14'b10100001101010;
9'd16   : cube_lut_4 = 14'b10100001101100;
9'd17   : cube_lut_4 = 14'b10100001101101;
9'd18   : cube_lut_4 = 14'b10100001101111;
9'd19   : cube_lut_4 = 14'b10100001110001;
9'd20   : cube_lut_4 = 14'b10100001110010;
9'd21   : cube_lut_4 = 14'b10100001110100;
9'd22   : cube_lut_4 = 14'b10100001110110;
9'd23   : cube_lut_4 = 14'b10100001110111;
9'd24   : cube_lut_4 = 14'b10100001111001;
9'd25   : cube_lut_4 = 14'b10100001111011;
9'd26   : cube_lut_4 = 14'b10100001111100;
9'd27   : cube_lut_4 = 14'b10100001111110;
9'd28   : cube_lut_4 = 14'b10100010000000;
9'd29   : cube_lut_4 = 14'b10100010000001;
9'd30   : cube_lut_4 = 14'b10100010000011;
9'd31   : cube_lut_4 = 14'b10100010000101;
9'd32   : cube_lut_4 = 14'b10100010000110;
9'd33   : cube_lut_4 = 14'b10100010001000;
9'd34   : cube_lut_4 = 14'b10100010001010;
9'd35   : cube_lut_4 = 14'b10100010001011;
9'd36   : cube_lut_4 = 14'b10100010001101;
9'd37   : cube_lut_4 = 14'b10100010001111;
9'd38   : cube_lut_4 = 14'b10100010010000;
9'd39   : cube_lut_4 = 14'b10100010010010;
9'd40   : cube_lut_4 = 14'b10100010010100;
9'd41   : cube_lut_4 = 14'b10100010010101;
9'd42   : cube_lut_4 = 14'b10100010010111;
9'd43   : cube_lut_4 = 14'b10100010011001;
9'd44   : cube_lut_4 = 14'b10100010011010;
9'd45   : cube_lut_4 = 14'b10100010011100;
9'd46   : cube_lut_4 = 14'b10100010011101;
9'd47   : cube_lut_4 = 14'b10100010011111;
9'd48   : cube_lut_4 = 14'b10100010100001;
9'd49   : cube_lut_4 = 14'b10100010100010;
9'd50   : cube_lut_4 = 14'b10100010100100;
9'd51   : cube_lut_4 = 14'b10100010100110;
9'd52   : cube_lut_4 = 14'b10100010100111;
9'd53   : cube_lut_4 = 14'b10100010101001;
9'd54   : cube_lut_4 = 14'b10100010101011;
9'd55   : cube_lut_4 = 14'b10100010101100;
9'd56   : cube_lut_4 = 14'b10100010101110;
9'd57   : cube_lut_4 = 14'b10100010110000;
9'd58   : cube_lut_4 = 14'b10100010110001;
9'd59   : cube_lut_4 = 14'b10100010110011;
9'd60   : cube_lut_4 = 14'b10100010110101;
9'd61   : cube_lut_4 = 14'b10100010110110;
9'd62   : cube_lut_4 = 14'b10100010111000;
9'd63   : cube_lut_4 = 14'b10100010111010;
9'd64   : cube_lut_4 = 14'b10100010111011;
9'd65   : cube_lut_4 = 14'b10100010111101;
9'd66   : cube_lut_4 = 14'b10100010111110;
9'd67   : cube_lut_4 = 14'b10100011000000;
9'd68   : cube_lut_4 = 14'b10100011000010;
9'd69   : cube_lut_4 = 14'b10100011000011;
9'd70   : cube_lut_4 = 14'b10100011000101;
9'd71   : cube_lut_4 = 14'b10100011000111;
9'd72   : cube_lut_4 = 14'b10100011001000;
9'd73   : cube_lut_4 = 14'b10100011001010;
9'd74   : cube_lut_4 = 14'b10100011001100;
9'd75   : cube_lut_4 = 14'b10100011001101;
9'd76   : cube_lut_4 = 14'b10100011001111;
9'd77   : cube_lut_4 = 14'b10100011010001;
9'd78   : cube_lut_4 = 14'b10100011010010;
9'd79   : cube_lut_4 = 14'b10100011010100;
9'd80   : cube_lut_4 = 14'b10100011010101;
9'd81   : cube_lut_4 = 14'b10100011010111;
9'd82   : cube_lut_4 = 14'b10100011011001;
9'd83   : cube_lut_4 = 14'b10100011011010;
9'd84   : cube_lut_4 = 14'b10100011011100;
9'd85   : cube_lut_4 = 14'b10100011011110;
9'd86   : cube_lut_4 = 14'b10100011011111;
9'd87   : cube_lut_4 = 14'b10100011100001;
9'd88   : cube_lut_4 = 14'b10100011100011;
9'd89   : cube_lut_4 = 14'b10100011100100;
9'd90   : cube_lut_4 = 14'b10100011100110;
9'd91   : cube_lut_4 = 14'b10100011100111;
9'd92   : cube_lut_4 = 14'b10100011101001;
9'd93   : cube_lut_4 = 14'b10100011101011;
9'd94   : cube_lut_4 = 14'b10100011101100;
9'd95   : cube_lut_4 = 14'b10100011101110;
9'd96   : cube_lut_4 = 14'b10100011110000;
9'd97   : cube_lut_4 = 14'b10100011110001;
9'd98   : cube_lut_4 = 14'b10100011110011;
9'd99   : cube_lut_4 = 14'b10100011110100;
9'd100   : cube_lut_4 = 14'b10100011110110;
9'd101   : cube_lut_4 = 14'b10100011111000;
9'd102   : cube_lut_4 = 14'b10100011111001;
9'd103   : cube_lut_4 = 14'b10100011111011;
9'd104   : cube_lut_4 = 14'b10100011111101;
9'd105   : cube_lut_4 = 14'b10100011111110;
9'd106   : cube_lut_4 = 14'b10100100000000;
9'd107   : cube_lut_4 = 14'b10100100000001;
9'd108   : cube_lut_4 = 14'b10100100000011;
9'd109   : cube_lut_4 = 14'b10100100000101;
9'd110   : cube_lut_4 = 14'b10100100000110;
9'd111   : cube_lut_4 = 14'b10100100001000;
9'd112   : cube_lut_4 = 14'b10100100001010;
9'd113   : cube_lut_4 = 14'b10100100001011;
9'd114   : cube_lut_4 = 14'b10100100001101;
9'd115   : cube_lut_4 = 14'b10100100001110;
9'd116   : cube_lut_4 = 14'b10100100010000;
9'd117   : cube_lut_4 = 14'b10100100010010;
9'd118   : cube_lut_4 = 14'b10100100010011;
9'd119   : cube_lut_4 = 14'b10100100010101;
9'd120   : cube_lut_4 = 14'b10100100010111;
9'd121   : cube_lut_4 = 14'b10100100011000;
9'd122   : cube_lut_4 = 14'b10100100011010;
9'd123   : cube_lut_4 = 14'b10100100011011;
9'd124   : cube_lut_4 = 14'b10100100011101;
9'd125   : cube_lut_4 = 14'b10100100011111;
9'd126   : cube_lut_4 = 14'b10100100100000;
9'd127   : cube_lut_4 = 14'b10100100100010;
9'd128   : cube_lut_4 = 14'b10100100100011;
9'd129   : cube_lut_4 = 14'b10100100100101;
9'd130   : cube_lut_4 = 14'b10100100100111;
9'd131   : cube_lut_4 = 14'b10100100101000;
9'd132   : cube_lut_4 = 14'b10100100101010;
9'd133   : cube_lut_4 = 14'b10100100101100;
9'd134   : cube_lut_4 = 14'b10100100101101;
9'd135   : cube_lut_4 = 14'b10100100101111;
9'd136   : cube_lut_4 = 14'b10100100110000;
9'd137   : cube_lut_4 = 14'b10100100110010;
9'd138   : cube_lut_4 = 14'b10100100110100;
9'd139   : cube_lut_4 = 14'b10100100110101;
9'd140   : cube_lut_4 = 14'b10100100110111;
9'd141   : cube_lut_4 = 14'b10100100111000;
9'd142   : cube_lut_4 = 14'b10100100111010;
9'd143   : cube_lut_4 = 14'b10100100111100;
9'd144   : cube_lut_4 = 14'b10100100111101;
9'd145   : cube_lut_4 = 14'b10100100111111;
9'd146   : cube_lut_4 = 14'b10100101000000;
9'd147   : cube_lut_4 = 14'b10100101000010;
9'd148   : cube_lut_4 = 14'b10100101000100;
9'd149   : cube_lut_4 = 14'b10100101000101;
9'd150   : cube_lut_4 = 14'b10100101000111;
9'd151   : cube_lut_4 = 14'b10100101001000;
9'd152   : cube_lut_4 = 14'b10100101001010;
9'd153   : cube_lut_4 = 14'b10100101001100;
9'd154   : cube_lut_4 = 14'b10100101001101;
9'd155   : cube_lut_4 = 14'b10100101001111;
9'd156   : cube_lut_4 = 14'b10100101010000;
9'd157   : cube_lut_4 = 14'b10100101010010;
9'd158   : cube_lut_4 = 14'b10100101010100;
9'd159   : cube_lut_4 = 14'b10100101010101;
9'd160   : cube_lut_4 = 14'b10100101010111;
9'd161   : cube_lut_4 = 14'b10100101011000;
9'd162   : cube_lut_4 = 14'b10100101011010;
9'd163   : cube_lut_4 = 14'b10100101011100;
9'd164   : cube_lut_4 = 14'b10100101011101;
9'd165   : cube_lut_4 = 14'b10100101011111;
9'd166   : cube_lut_4 = 14'b10100101100000;
9'd167   : cube_lut_4 = 14'b10100101100010;
9'd168   : cube_lut_4 = 14'b10100101100100;
9'd169   : cube_lut_4 = 14'b10100101100101;
9'd170   : cube_lut_4 = 14'b10100101100111;
9'd171   : cube_lut_4 = 14'b10100101101000;
9'd172   : cube_lut_4 = 14'b10100101101010;
9'd173   : cube_lut_4 = 14'b10100101101100;
9'd174   : cube_lut_4 = 14'b10100101101101;
9'd175   : cube_lut_4 = 14'b10100101101111;
9'd176   : cube_lut_4 = 14'b10100101110000;
9'd177   : cube_lut_4 = 14'b10100101110010;
9'd178   : cube_lut_4 = 14'b10100101110100;
9'd179   : cube_lut_4 = 14'b10100101110101;
9'd180   : cube_lut_4 = 14'b10100101110111;
9'd181   : cube_lut_4 = 14'b10100101111000;
9'd182   : cube_lut_4 = 14'b10100101111010;
9'd183   : cube_lut_4 = 14'b10100101111011;
9'd184   : cube_lut_4 = 14'b10100101111101;
9'd185   : cube_lut_4 = 14'b10100101111111;
9'd186   : cube_lut_4 = 14'b10100110000000;
9'd187   : cube_lut_4 = 14'b10100110000010;
9'd188   : cube_lut_4 = 14'b10100110000011;
9'd189   : cube_lut_4 = 14'b10100110000101;
9'd190   : cube_lut_4 = 14'b10100110000111;
9'd191   : cube_lut_4 = 14'b10100110001000;
9'd192   : cube_lut_4 = 14'b10100110001010;
9'd193   : cube_lut_4 = 14'b10100110001011;
9'd194   : cube_lut_4 = 14'b10100110001101;
9'd195   : cube_lut_4 = 14'b10100110001110;
9'd196   : cube_lut_4 = 14'b10100110010000;
9'd197   : cube_lut_4 = 14'b10100110010010;
9'd198   : cube_lut_4 = 14'b10100110010011;
9'd199   : cube_lut_4 = 14'b10100110010101;
9'd200   : cube_lut_4 = 14'b10100110010110;
9'd201   : cube_lut_4 = 14'b10100110011000;
9'd202   : cube_lut_4 = 14'b10100110011010;
9'd203   : cube_lut_4 = 14'b10100110011011;
9'd204   : cube_lut_4 = 14'b10100110011101;
9'd205   : cube_lut_4 = 14'b10100110011110;
9'd206   : cube_lut_4 = 14'b10100110100000;
9'd207   : cube_lut_4 = 14'b10100110100001;
9'd208   : cube_lut_4 = 14'b10100110100011;
9'd209   : cube_lut_4 = 14'b10100110100101;
9'd210   : cube_lut_4 = 14'b10100110100110;
9'd211   : cube_lut_4 = 14'b10100110101000;
9'd212   : cube_lut_4 = 14'b10100110101001;
9'd213   : cube_lut_4 = 14'b10100110101011;
9'd214   : cube_lut_4 = 14'b10100110101100;
9'd215   : cube_lut_4 = 14'b10100110101110;
9'd216   : cube_lut_4 = 14'b10100110110000;
9'd217   : cube_lut_4 = 14'b10100110110001;
9'd218   : cube_lut_4 = 14'b10100110110011;
9'd219   : cube_lut_4 = 14'b10100110110100;
9'd220   : cube_lut_4 = 14'b10100110110110;
9'd221   : cube_lut_4 = 14'b10100110110111;
9'd222   : cube_lut_4 = 14'b10100110111001;
9'd223   : cube_lut_4 = 14'b10100110111011;
9'd224   : cube_lut_4 = 14'b10100110111100;
9'd225   : cube_lut_4 = 14'b10100110111110;
9'd226   : cube_lut_4 = 14'b10100110111111;
9'd227   : cube_lut_4 = 14'b10100111000001;
9'd228   : cube_lut_4 = 14'b10100111000010;
9'd229   : cube_lut_4 = 14'b10100111000100;
9'd230   : cube_lut_4 = 14'b10100111000110;
9'd231   : cube_lut_4 = 14'b10100111000111;
9'd232   : cube_lut_4 = 14'b10100111001001;
9'd233   : cube_lut_4 = 14'b10100111001010;
9'd234   : cube_lut_4 = 14'b10100111001100;
9'd235   : cube_lut_4 = 14'b10100111001101;
9'd236   : cube_lut_4 = 14'b10100111001111;
9'd237   : cube_lut_4 = 14'b10100111010000;
9'd238   : cube_lut_4 = 14'b10100111010010;
9'd239   : cube_lut_4 = 14'b10100111010100;
9'd240   : cube_lut_4 = 14'b10100111010101;
9'd241   : cube_lut_4 = 14'b10100111010111;
9'd242   : cube_lut_4 = 14'b10100111011000;
9'd243   : cube_lut_4 = 14'b10100111011010;
9'd244   : cube_lut_4 = 14'b10100111011011;
9'd245   : cube_lut_4 = 14'b10100111011101;
9'd246   : cube_lut_4 = 14'b10100111011111;
9'd247   : cube_lut_4 = 14'b10100111100000;
9'd248   : cube_lut_4 = 14'b10100111100010;
9'd249   : cube_lut_4 = 14'b10100111100011;
9'd250   : cube_lut_4 = 14'b10100111100101;
9'd251   : cube_lut_4 = 14'b10100111100110;
9'd252   : cube_lut_4 = 14'b10100111101000;
9'd253   : cube_lut_4 = 14'b10100111101001;
9'd254   : cube_lut_4 = 14'b10100111101011;
9'd255   : cube_lut_4 = 14'b10100111101101;
9'd256   : cube_lut_4 = 14'b10100111101110;
9'd257   : cube_lut_4 = 14'b10100111110000;
9'd258   : cube_lut_4 = 14'b10100111110001;
9'd259   : cube_lut_4 = 14'b10100111110011;
9'd260   : cube_lut_4 = 14'b10100111110100;
9'd261   : cube_lut_4 = 14'b10100111110110;
9'd262   : cube_lut_4 = 14'b10100111110111;
9'd263   : cube_lut_4 = 14'b10100111111001;
9'd264   : cube_lut_4 = 14'b10100111111010;
9'd265   : cube_lut_4 = 14'b10100111111100;
9'd266   : cube_lut_4 = 14'b10100111111110;
9'd267   : cube_lut_4 = 14'b10100111111111;
9'd268   : cube_lut_4 = 14'b10101000000001;
9'd269   : cube_lut_4 = 14'b10101000000010;
9'd270   : cube_lut_4 = 14'b10101000000100;
9'd271   : cube_lut_4 = 14'b10101000000101;
9'd272   : cube_lut_4 = 14'b10101000000111;
9'd273   : cube_lut_4 = 14'b10101000001000;
9'd274   : cube_lut_4 = 14'b10101000001010;
9'd275   : cube_lut_4 = 14'b10101000001011;
9'd276   : cube_lut_4 = 14'b10101000001101;
9'd277   : cube_lut_4 = 14'b10101000001111;
9'd278   : cube_lut_4 = 14'b10101000010000;
9'd279   : cube_lut_4 = 14'b10101000010010;
9'd280   : cube_lut_4 = 14'b10101000010011;
9'd281   : cube_lut_4 = 14'b10101000010101;
9'd282   : cube_lut_4 = 14'b10101000010110;
9'd283   : cube_lut_4 = 14'b10101000011000;
9'd284   : cube_lut_4 = 14'b10101000011001;
9'd285   : cube_lut_4 = 14'b10101000011011;
9'd286   : cube_lut_4 = 14'b10101000011100;
9'd287   : cube_lut_4 = 14'b10101000011110;
9'd288   : cube_lut_4 = 14'b10101000100000;
9'd289   : cube_lut_4 = 14'b10101000100001;
9'd290   : cube_lut_4 = 14'b10101000100011;
9'd291   : cube_lut_4 = 14'b10101000100100;
9'd292   : cube_lut_4 = 14'b10101000100110;
9'd293   : cube_lut_4 = 14'b10101000100111;
9'd294   : cube_lut_4 = 14'b10101000101001;
9'd295   : cube_lut_4 = 14'b10101000101010;
9'd296   : cube_lut_4 = 14'b10101000101100;
9'd297   : cube_lut_4 = 14'b10101000101101;
9'd298   : cube_lut_4 = 14'b10101000101111;
9'd299   : cube_lut_4 = 14'b10101000110000;
9'd300   : cube_lut_4 = 14'b10101000110010;
9'd301   : cube_lut_4 = 14'b10101000110011;
9'd302   : cube_lut_4 = 14'b10101000110101;
9'd303   : cube_lut_4 = 14'b10101000110111;
9'd304   : cube_lut_4 = 14'b10101000111000;
9'd305   : cube_lut_4 = 14'b10101000111010;
9'd306   : cube_lut_4 = 14'b10101000111011;
9'd307   : cube_lut_4 = 14'b10101000111101;
9'd308   : cube_lut_4 = 14'b10101000111110;
9'd309   : cube_lut_4 = 14'b10101001000000;
9'd310   : cube_lut_4 = 14'b10101001000001;
9'd311   : cube_lut_4 = 14'b10101001000011;
9'd312   : cube_lut_4 = 14'b10101001000100;
9'd313   : cube_lut_4 = 14'b10101001000110;
9'd314   : cube_lut_4 = 14'b10101001000111;
9'd315   : cube_lut_4 = 14'b10101001001001;
9'd316   : cube_lut_4 = 14'b10101001001010;
9'd317   : cube_lut_4 = 14'b10101001001100;
9'd318   : cube_lut_4 = 14'b10101001001101;
9'd319   : cube_lut_4 = 14'b10101001001111;
9'd320   : cube_lut_4 = 14'b10101001010001;
9'd321   : cube_lut_4 = 14'b10101001010010;
9'd322   : cube_lut_4 = 14'b10101001010100;
9'd323   : cube_lut_4 = 14'b10101001010101;
9'd324   : cube_lut_4 = 14'b10101001010111;
9'd325   : cube_lut_4 = 14'b10101001011000;
9'd326   : cube_lut_4 = 14'b10101001011010;
9'd327   : cube_lut_4 = 14'b10101001011011;
9'd328   : cube_lut_4 = 14'b10101001011101;
9'd329   : cube_lut_4 = 14'b10101001011110;
9'd330   : cube_lut_4 = 14'b10101001100000;
9'd331   : cube_lut_4 = 14'b10101001100001;
9'd332   : cube_lut_4 = 14'b10101001100011;
9'd333   : cube_lut_4 = 14'b10101001100100;
9'd334   : cube_lut_4 = 14'b10101001100110;
9'd335   : cube_lut_4 = 14'b10101001100111;
9'd336   : cube_lut_4 = 14'b10101001101001;
9'd337   : cube_lut_4 = 14'b10101001101010;
9'd338   : cube_lut_4 = 14'b10101001101100;
9'd339   : cube_lut_4 = 14'b10101001101101;
9'd340   : cube_lut_4 = 14'b10101001101111;
9'd341   : cube_lut_4 = 14'b10101001110000;
9'd342   : cube_lut_4 = 14'b10101001110010;
9'd343   : cube_lut_4 = 14'b10101001110100;
9'd344   : cube_lut_4 = 14'b10101001110101;
9'd345   : cube_lut_4 = 14'b10101001110111;
9'd346   : cube_lut_4 = 14'b10101001111000;
9'd347   : cube_lut_4 = 14'b10101001111010;
9'd348   : cube_lut_4 = 14'b10101001111011;
9'd349   : cube_lut_4 = 14'b10101001111101;
9'd350   : cube_lut_4 = 14'b10101001111110;
9'd351   : cube_lut_4 = 14'b10101010000000;
9'd352   : cube_lut_4 = 14'b10101010000001;
9'd353   : cube_lut_4 = 14'b10101010000011;
9'd354   : cube_lut_4 = 14'b10101010000100;
9'd355   : cube_lut_4 = 14'b10101010000110;
9'd356   : cube_lut_4 = 14'b10101010000111;
9'd357   : cube_lut_4 = 14'b10101010001001;
9'd358   : cube_lut_4 = 14'b10101010001010;
9'd359   : cube_lut_4 = 14'b10101010001100;
9'd360   : cube_lut_4 = 14'b10101010001101;
9'd361   : cube_lut_4 = 14'b10101010001111;
9'd362   : cube_lut_4 = 14'b10101010010000;
9'd363   : cube_lut_4 = 14'b10101010010010;
9'd364   : cube_lut_4 = 14'b10101010010011;
9'd365   : cube_lut_4 = 14'b10101010010101;
9'd366   : cube_lut_4 = 14'b10101010010110;
9'd367   : cube_lut_4 = 14'b10101010011000;
9'd368   : cube_lut_4 = 14'b10101010011001;
9'd369   : cube_lut_4 = 14'b10101010011011;
9'd370   : cube_lut_4 = 14'b10101010011100;
9'd371   : cube_lut_4 = 14'b10101010011110;
9'd372   : cube_lut_4 = 14'b10101010011111;
9'd373   : cube_lut_4 = 14'b10101010100001;
9'd374   : cube_lut_4 = 14'b10101010100010;
9'd375   : cube_lut_4 = 14'b10101010100100;
9'd376   : cube_lut_4 = 14'b10101010100101;
9'd377   : cube_lut_4 = 14'b10101010100111;
9'd378   : cube_lut_4 = 14'b10101010101000;
9'd379   : cube_lut_4 = 14'b10101010101010;
9'd380   : cube_lut_4 = 14'b10101010101011;
9'd381   : cube_lut_4 = 14'b10101010101101;
9'd382   : cube_lut_4 = 14'b10101010101110;
9'd383   : cube_lut_4 = 14'b10101010110000;
9'd384   : cube_lut_4 = 14'b10101010110001;
9'd385   : cube_lut_4 = 14'b10101010110011;
9'd386   : cube_lut_4 = 14'b10101010110100;
9'd387   : cube_lut_4 = 14'b10101010110110;
9'd388   : cube_lut_4 = 14'b10101010110111;
9'd389   : cube_lut_4 = 14'b10101010111001;
9'd390   : cube_lut_4 = 14'b10101010111010;
9'd391   : cube_lut_4 = 14'b10101010111100;
9'd392   : cube_lut_4 = 14'b10101010111101;
9'd393   : cube_lut_4 = 14'b10101010111111;
9'd394   : cube_lut_4 = 14'b10101011000000;
9'd395   : cube_lut_4 = 14'b10101011000010;
9'd396   : cube_lut_4 = 14'b10101011000011;
9'd397   : cube_lut_4 = 14'b10101011000101;
9'd398   : cube_lut_4 = 14'b10101011000110;
9'd399   : cube_lut_4 = 14'b10101011001000;
9'd400   : cube_lut_4 = 14'b10101011001001;
9'd401   : cube_lut_4 = 14'b10101011001011;
9'd402   : cube_lut_4 = 14'b10101011001100;
9'd403   : cube_lut_4 = 14'b10101011001110;
9'd404   : cube_lut_4 = 14'b10101011001111;
9'd405   : cube_lut_4 = 14'b10101011010001;
9'd406   : cube_lut_4 = 14'b10101011010010;
9'd407   : cube_lut_4 = 14'b10101011010100;
9'd408   : cube_lut_4 = 14'b10101011010101;
9'd409   : cube_lut_4 = 14'b10101011010111;
9'd410   : cube_lut_4 = 14'b10101011011000;
9'd411   : cube_lut_4 = 14'b10101011011010;
9'd412   : cube_lut_4 = 14'b10101011011011;
9'd413   : cube_lut_4 = 14'b10101011011101;
9'd414   : cube_lut_4 = 14'b10101011011110;
9'd415   : cube_lut_4 = 14'b10101011100000;
9'd416   : cube_lut_4 = 14'b10101011100001;
9'd417   : cube_lut_4 = 14'b10101011100010;
9'd418   : cube_lut_4 = 14'b10101011100100;
9'd419   : cube_lut_4 = 14'b10101011100101;
9'd420   : cube_lut_4 = 14'b10101011100111;
9'd421   : cube_lut_4 = 14'b10101011101000;
9'd422   : cube_lut_4 = 14'b10101011101010;
9'd423   : cube_lut_4 = 14'b10101011101011;
9'd424   : cube_lut_4 = 14'b10101011101101;
9'd425   : cube_lut_4 = 14'b10101011101110;
9'd426   : cube_lut_4 = 14'b10101011110000;
9'd427   : cube_lut_4 = 14'b10101011110001;
9'd428   : cube_lut_4 = 14'b10101011110011;
9'd429   : cube_lut_4 = 14'b10101011110100;
9'd430   : cube_lut_4 = 14'b10101011110110;
9'd431   : cube_lut_4 = 14'b10101011110111;
9'd432   : cube_lut_4 = 14'b10101011111001;
9'd433   : cube_lut_4 = 14'b10101011111010;
9'd434   : cube_lut_4 = 14'b10101011111100;
9'd435   : cube_lut_4 = 14'b10101011111101;
9'd436   : cube_lut_4 = 14'b10101011111111;
9'd437   : cube_lut_4 = 14'b10101100000000;
9'd438   : cube_lut_4 = 14'b10101100000010;
9'd439   : cube_lut_4 = 14'b10101100000011;
9'd440   : cube_lut_4 = 14'b10101100000101;
9'd441   : cube_lut_4 = 14'b10101100000110;
9'd442   : cube_lut_4 = 14'b10101100000111;
9'd443   : cube_lut_4 = 14'b10101100001001;
9'd444   : cube_lut_4 = 14'b10101100001010;
9'd445   : cube_lut_4 = 14'b10101100001100;
9'd446   : cube_lut_4 = 14'b10101100001101;
9'd447   : cube_lut_4 = 14'b10101100001111;
9'd448   : cube_lut_4 = 14'b10101100010000;
9'd449   : cube_lut_4 = 14'b10101100010010;
9'd450   : cube_lut_4 = 14'b10101100010011;
9'd451   : cube_lut_4 = 14'b10101100010101;
9'd452   : cube_lut_4 = 14'b10101100010110;
9'd453   : cube_lut_4 = 14'b10101100011000;
9'd454   : cube_lut_4 = 14'b10101100011001;
9'd455   : cube_lut_4 = 14'b10101100011011;
9'd456   : cube_lut_4 = 14'b10101100011100;
9'd457   : cube_lut_4 = 14'b10101100011110;
9'd458   : cube_lut_4 = 14'b10101100011111;
9'd459   : cube_lut_4 = 14'b10101100100000;
9'd460   : cube_lut_4 = 14'b10101100100010;
9'd461   : cube_lut_4 = 14'b10101100100011;
9'd462   : cube_lut_4 = 14'b10101100100101;
9'd463   : cube_lut_4 = 14'b10101100100110;
9'd464   : cube_lut_4 = 14'b10101100101000;
9'd465   : cube_lut_4 = 14'b10101100101001;
9'd466   : cube_lut_4 = 14'b10101100101011;
9'd467   : cube_lut_4 = 14'b10101100101100;
9'd468   : cube_lut_4 = 14'b10101100101110;
9'd469   : cube_lut_4 = 14'b10101100101111;
9'd470   : cube_lut_4 = 14'b10101100110001;
9'd471   : cube_lut_4 = 14'b10101100110010;
9'd472   : cube_lut_4 = 14'b10101100110100;
9'd473   : cube_lut_4 = 14'b10101100110101;
9'd474   : cube_lut_4 = 14'b10101100110110;
9'd475   : cube_lut_4 = 14'b10101100111000;
9'd476   : cube_lut_4 = 14'b10101100111001;
9'd477   : cube_lut_4 = 14'b10101100111011;
9'd478   : cube_lut_4 = 14'b10101100111100;
9'd479   : cube_lut_4 = 14'b10101100111110;
9'd480   : cube_lut_4 = 14'b10101100111111;
9'd481   : cube_lut_4 = 14'b10101101000001;
9'd482   : cube_lut_4 = 14'b10101101000010;
9'd483   : cube_lut_4 = 14'b10101101000100;
9'd484   : cube_lut_4 = 14'b10101101000101;
9'd485   : cube_lut_4 = 14'b10101101000111;
9'd486   : cube_lut_4 = 14'b10101101001000;
9'd487   : cube_lut_4 = 14'b10101101001001;
9'd488   : cube_lut_4 = 14'b10101101001011;
9'd489   : cube_lut_4 = 14'b10101101001100;
9'd490   : cube_lut_4 = 14'b10101101001110;
9'd491   : cube_lut_4 = 14'b10101101001111;
9'd492   : cube_lut_4 = 14'b10101101010001;
9'd493   : cube_lut_4 = 14'b10101101010010;
9'd494   : cube_lut_4 = 14'b10101101010100;
9'd495   : cube_lut_4 = 14'b10101101010101;
9'd496   : cube_lut_4 = 14'b10101101010111;
9'd497   : cube_lut_4 = 14'b10101101011000;
9'd498   : cube_lut_4 = 14'b10101101011001;
9'd499   : cube_lut_4 = 14'b10101101011011;
9'd500   : cube_lut_4 = 14'b10101101011100;
9'd501   : cube_lut_4 = 14'b10101101011110;
9'd502   : cube_lut_4 = 14'b10101101011111;
9'd503   : cube_lut_4 = 14'b10101101100001;
9'd504   : cube_lut_4 = 14'b10101101100010;
9'd505   : cube_lut_4 = 14'b10101101100100;
9'd506   : cube_lut_4 = 14'b10101101100101;
9'd507   : cube_lut_4 = 14'b10101101100111;
9'd508   : cube_lut_4 = 14'b10101101101000;
9'd509   : cube_lut_4 = 14'b10101101101001;
9'd510   : cube_lut_4 = 14'b10101101101011;
9'd511   : cube_lut_4 = 14'b10101101101100;

    endcase
end

always@* begin
    
    cube_lut_5 = 0;
    
    case(i_data[8:0])
 
 9'd0   : cube_lut_5 = 14'b10101101101110;
9'd1   : cube_lut_5 = 14'b10101101101111;
9'd2   : cube_lut_5 = 14'b10101101110001;
9'd3   : cube_lut_5 = 14'b10101101110010;
9'd4   : cube_lut_5 = 14'b10101101110100;
9'd5   : cube_lut_5 = 14'b10101101110101;
9'd6   : cube_lut_5 = 14'b10101101110110;
9'd7   : cube_lut_5 = 14'b10101101111000;
9'd8   : cube_lut_5 = 14'b10101101111001;
9'd9   : cube_lut_5 = 14'b10101101111011;
9'd10   : cube_lut_5 = 14'b10101101111100;
9'd11   : cube_lut_5 = 14'b10101101111110;
9'd12   : cube_lut_5 = 14'b10101101111111;
9'd13   : cube_lut_5 = 14'b10101110000001;
9'd14   : cube_lut_5 = 14'b10101110000010;
9'd15   : cube_lut_5 = 14'b10101110000011;
9'd16   : cube_lut_5 = 14'b10101110000101;
9'd17   : cube_lut_5 = 14'b10101110000110;
9'd18   : cube_lut_5 = 14'b10101110001000;
9'd19   : cube_lut_5 = 14'b10101110001001;
9'd20   : cube_lut_5 = 14'b10101110001011;
9'd21   : cube_lut_5 = 14'b10101110001100;
9'd22   : cube_lut_5 = 14'b10101110001110;
9'd23   : cube_lut_5 = 14'b10101110001111;
9'd24   : cube_lut_5 = 14'b10101110010000;
9'd25   : cube_lut_5 = 14'b10101110010010;
9'd26   : cube_lut_5 = 14'b10101110010011;
9'd27   : cube_lut_5 = 14'b10101110010101;
9'd28   : cube_lut_5 = 14'b10101110010110;
9'd29   : cube_lut_5 = 14'b10101110011000;
9'd30   : cube_lut_5 = 14'b10101110011001;
9'd31   : cube_lut_5 = 14'b10101110011010;
9'd32   : cube_lut_5 = 14'b10101110011100;
9'd33   : cube_lut_5 = 14'b10101110011101;
9'd34   : cube_lut_5 = 14'b10101110011111;
9'd35   : cube_lut_5 = 14'b10101110100000;
9'd36   : cube_lut_5 = 14'b10101110100010;
9'd37   : cube_lut_5 = 14'b10101110100011;
9'd38   : cube_lut_5 = 14'b10101110100100;
9'd39   : cube_lut_5 = 14'b10101110100110;
9'd40   : cube_lut_5 = 14'b10101110100111;
9'd41   : cube_lut_5 = 14'b10101110101001;
9'd42   : cube_lut_5 = 14'b10101110101010;
9'd43   : cube_lut_5 = 14'b10101110101100;
9'd44   : cube_lut_5 = 14'b10101110101101;
9'd45   : cube_lut_5 = 14'b10101110101111;
9'd46   : cube_lut_5 = 14'b10101110110000;
9'd47   : cube_lut_5 = 14'b10101110110001;
9'd48   : cube_lut_5 = 14'b10101110110011;
9'd49   : cube_lut_5 = 14'b10101110110100;
9'd50   : cube_lut_5 = 14'b10101110110110;
9'd51   : cube_lut_5 = 14'b10101110110111;
9'd52   : cube_lut_5 = 14'b10101110111001;
9'd53   : cube_lut_5 = 14'b10101110111010;
9'd54   : cube_lut_5 = 14'b10101110111011;
9'd55   : cube_lut_5 = 14'b10101110111101;
9'd56   : cube_lut_5 = 14'b10101110111110;
9'd57   : cube_lut_5 = 14'b10101111000000;
9'd58   : cube_lut_5 = 14'b10101111000001;
9'd59   : cube_lut_5 = 14'b10101111000011;
9'd60   : cube_lut_5 = 14'b10101111000100;
9'd61   : cube_lut_5 = 14'b10101111000101;
9'd62   : cube_lut_5 = 14'b10101111000111;
9'd63   : cube_lut_5 = 14'b10101111001000;
9'd64   : cube_lut_5 = 14'b10101111001010;
9'd65   : cube_lut_5 = 14'b10101111001011;
9'd66   : cube_lut_5 = 14'b10101111001100;
9'd67   : cube_lut_5 = 14'b10101111001110;
9'd68   : cube_lut_5 = 14'b10101111001111;
9'd69   : cube_lut_5 = 14'b10101111010001;
9'd70   : cube_lut_5 = 14'b10101111010010;
9'd71   : cube_lut_5 = 14'b10101111010100;
9'd72   : cube_lut_5 = 14'b10101111010101;
9'd73   : cube_lut_5 = 14'b10101111010110;
9'd74   : cube_lut_5 = 14'b10101111011000;
9'd75   : cube_lut_5 = 14'b10101111011001;
9'd76   : cube_lut_5 = 14'b10101111011011;
9'd77   : cube_lut_5 = 14'b10101111011100;
9'd78   : cube_lut_5 = 14'b10101111011110;
9'd79   : cube_lut_5 = 14'b10101111011111;
9'd80   : cube_lut_5 = 14'b10101111100000;
9'd81   : cube_lut_5 = 14'b10101111100010;
9'd82   : cube_lut_5 = 14'b10101111100011;
9'd83   : cube_lut_5 = 14'b10101111100101;
9'd84   : cube_lut_5 = 14'b10101111100110;
9'd85   : cube_lut_5 = 14'b10101111100111;
9'd86   : cube_lut_5 = 14'b10101111101001;
9'd87   : cube_lut_5 = 14'b10101111101010;
9'd88   : cube_lut_5 = 14'b10101111101100;
9'd89   : cube_lut_5 = 14'b10101111101101;
9'd90   : cube_lut_5 = 14'b10101111101111;
9'd91   : cube_lut_5 = 14'b10101111110000;
9'd92   : cube_lut_5 = 14'b10101111110001;
9'd93   : cube_lut_5 = 14'b10101111110011;
9'd94   : cube_lut_5 = 14'b10101111110100;
9'd95   : cube_lut_5 = 14'b10101111110110;
9'd96   : cube_lut_5 = 14'b10101111110111;
9'd97   : cube_lut_5 = 14'b10101111111000;
9'd98   : cube_lut_5 = 14'b10101111111010;
9'd99   : cube_lut_5 = 14'b10101111111011;
9'd100   : cube_lut_5 = 14'b10101111111101;
9'd101   : cube_lut_5 = 14'b10101111111110;
9'd102   : cube_lut_5 = 14'b10110000000000;
9'd103   : cube_lut_5 = 14'b10110000000001;
9'd104   : cube_lut_5 = 14'b10110000000010;
9'd105   : cube_lut_5 = 14'b10110000000100;
9'd106   : cube_lut_5 = 14'b10110000000101;
9'd107   : cube_lut_5 = 14'b10110000000111;
9'd108   : cube_lut_5 = 14'b10110000001000;
9'd109   : cube_lut_5 = 14'b10110000001001;
9'd110   : cube_lut_5 = 14'b10110000001011;
9'd111   : cube_lut_5 = 14'b10110000001100;
9'd112   : cube_lut_5 = 14'b10110000001110;
9'd113   : cube_lut_5 = 14'b10110000001111;
9'd114   : cube_lut_5 = 14'b10110000010000;
9'd115   : cube_lut_5 = 14'b10110000010010;
9'd116   : cube_lut_5 = 14'b10110000010011;
9'd117   : cube_lut_5 = 14'b10110000010101;
9'd118   : cube_lut_5 = 14'b10110000010110;
9'd119   : cube_lut_5 = 14'b10110000010111;
9'd120   : cube_lut_5 = 14'b10110000011001;
9'd121   : cube_lut_5 = 14'b10110000011010;
9'd122   : cube_lut_5 = 14'b10110000011100;
9'd123   : cube_lut_5 = 14'b10110000011101;
9'd124   : cube_lut_5 = 14'b10110000011110;
9'd125   : cube_lut_5 = 14'b10110000100000;
9'd126   : cube_lut_5 = 14'b10110000100001;
9'd127   : cube_lut_5 = 14'b10110000100011;
9'd128   : cube_lut_5 = 14'b10110000100100;
9'd129   : cube_lut_5 = 14'b10110000100101;
9'd130   : cube_lut_5 = 14'b10110000100111;
9'd131   : cube_lut_5 = 14'b10110000101000;
9'd132   : cube_lut_5 = 14'b10110000101010;
9'd133   : cube_lut_5 = 14'b10110000101011;
9'd134   : cube_lut_5 = 14'b10110000101100;
9'd135   : cube_lut_5 = 14'b10110000101110;
9'd136   : cube_lut_5 = 14'b10110000101111;
9'd137   : cube_lut_5 = 14'b10110000110001;
9'd138   : cube_lut_5 = 14'b10110000110010;
9'd139   : cube_lut_5 = 14'b10110000110011;
9'd140   : cube_lut_5 = 14'b10110000110101;
9'd141   : cube_lut_5 = 14'b10110000110110;
9'd142   : cube_lut_5 = 14'b10110000111000;
9'd143   : cube_lut_5 = 14'b10110000111001;
9'd144   : cube_lut_5 = 14'b10110000111010;
9'd145   : cube_lut_5 = 14'b10110000111100;
9'd146   : cube_lut_5 = 14'b10110000111101;
9'd147   : cube_lut_5 = 14'b10110000111111;
9'd148   : cube_lut_5 = 14'b10110001000000;
9'd149   : cube_lut_5 = 14'b10110001000001;
9'd150   : cube_lut_5 = 14'b10110001000011;
9'd151   : cube_lut_5 = 14'b10110001000100;
9'd152   : cube_lut_5 = 14'b10110001000110;
9'd153   : cube_lut_5 = 14'b10110001000111;
9'd154   : cube_lut_5 = 14'b10110001001000;
9'd155   : cube_lut_5 = 14'b10110001001010;
9'd156   : cube_lut_5 = 14'b10110001001011;
9'd157   : cube_lut_5 = 14'b10110001001101;
9'd158   : cube_lut_5 = 14'b10110001001110;
9'd159   : cube_lut_5 = 14'b10110001001111;
9'd160   : cube_lut_5 = 14'b10110001010001;
9'd161   : cube_lut_5 = 14'b10110001010010;
9'd162   : cube_lut_5 = 14'b10110001010100;
9'd163   : cube_lut_5 = 14'b10110001010101;
9'd164   : cube_lut_5 = 14'b10110001010110;
9'd165   : cube_lut_5 = 14'b10110001011000;
9'd166   : cube_lut_5 = 14'b10110001011001;
9'd167   : cube_lut_5 = 14'b10110001011010;
9'd168   : cube_lut_5 = 14'b10110001011100;
9'd169   : cube_lut_5 = 14'b10110001011101;
9'd170   : cube_lut_5 = 14'b10110001011111;
9'd171   : cube_lut_5 = 14'b10110001100000;
9'd172   : cube_lut_5 = 14'b10110001100001;
9'd173   : cube_lut_5 = 14'b10110001100011;
9'd174   : cube_lut_5 = 14'b10110001100100;
9'd175   : cube_lut_5 = 14'b10110001100110;
9'd176   : cube_lut_5 = 14'b10110001100111;
9'd177   : cube_lut_5 = 14'b10110001101000;
9'd178   : cube_lut_5 = 14'b10110001101010;
9'd179   : cube_lut_5 = 14'b10110001101011;
9'd180   : cube_lut_5 = 14'b10110001101100;
9'd181   : cube_lut_5 = 14'b10110001101110;
9'd182   : cube_lut_5 = 14'b10110001101111;
9'd183   : cube_lut_5 = 14'b10110001110001;
9'd184   : cube_lut_5 = 14'b10110001110010;
9'd185   : cube_lut_5 = 14'b10110001110011;
9'd186   : cube_lut_5 = 14'b10110001110101;
9'd187   : cube_lut_5 = 14'b10110001110110;
9'd188   : cube_lut_5 = 14'b10110001111000;
9'd189   : cube_lut_5 = 14'b10110001111001;
9'd190   : cube_lut_5 = 14'b10110001111010;
9'd191   : cube_lut_5 = 14'b10110001111100;
9'd192   : cube_lut_5 = 14'b10110001111101;
9'd193   : cube_lut_5 = 14'b10110001111110;
9'd194   : cube_lut_5 = 14'b10110010000000;
9'd195   : cube_lut_5 = 14'b10110010000001;
9'd196   : cube_lut_5 = 14'b10110010000011;
9'd197   : cube_lut_5 = 14'b10110010000100;
9'd198   : cube_lut_5 = 14'b10110010000101;
9'd199   : cube_lut_5 = 14'b10110010000111;
9'd200   : cube_lut_5 = 14'b10110010001000;
9'd201   : cube_lut_5 = 14'b10110010001001;
9'd202   : cube_lut_5 = 14'b10110010001011;
9'd203   : cube_lut_5 = 14'b10110010001100;
9'd204   : cube_lut_5 = 14'b10110010001110;
9'd205   : cube_lut_5 = 14'b10110010001111;
9'd206   : cube_lut_5 = 14'b10110010010000;
9'd207   : cube_lut_5 = 14'b10110010010010;
9'd208   : cube_lut_5 = 14'b10110010010011;
9'd209   : cube_lut_5 = 14'b10110010010100;
9'd210   : cube_lut_5 = 14'b10110010010110;
9'd211   : cube_lut_5 = 14'b10110010010111;
9'd212   : cube_lut_5 = 14'b10110010011001;
9'd213   : cube_lut_5 = 14'b10110010011010;
9'd214   : cube_lut_5 = 14'b10110010011011;
9'd215   : cube_lut_5 = 14'b10110010011101;
9'd216   : cube_lut_5 = 14'b10110010011110;
9'd217   : cube_lut_5 = 14'b10110010011111;
9'd218   : cube_lut_5 = 14'b10110010100001;
9'd219   : cube_lut_5 = 14'b10110010100010;
9'd220   : cube_lut_5 = 14'b10110010100100;
9'd221   : cube_lut_5 = 14'b10110010100101;
9'd222   : cube_lut_5 = 14'b10110010100110;
9'd223   : cube_lut_5 = 14'b10110010101000;
9'd224   : cube_lut_5 = 14'b10110010101001;
9'd225   : cube_lut_5 = 14'b10110010101010;
9'd226   : cube_lut_5 = 14'b10110010101100;
9'd227   : cube_lut_5 = 14'b10110010101101;
9'd228   : cube_lut_5 = 14'b10110010101110;
9'd229   : cube_lut_5 = 14'b10110010110000;
9'd230   : cube_lut_5 = 14'b10110010110001;
9'd231   : cube_lut_5 = 14'b10110010110011;
9'd232   : cube_lut_5 = 14'b10110010110100;
9'd233   : cube_lut_5 = 14'b10110010110101;
9'd234   : cube_lut_5 = 14'b10110010110111;
9'd235   : cube_lut_5 = 14'b10110010111000;
9'd236   : cube_lut_5 = 14'b10110010111001;
9'd237   : cube_lut_5 = 14'b10110010111011;
9'd238   : cube_lut_5 = 14'b10110010111100;
9'd239   : cube_lut_5 = 14'b10110010111110;
9'd240   : cube_lut_5 = 14'b10110010111111;
9'd241   : cube_lut_5 = 14'b10110011000000;
9'd242   : cube_lut_5 = 14'b10110011000010;
9'd243   : cube_lut_5 = 14'b10110011000011;
9'd244   : cube_lut_5 = 14'b10110011000100;
9'd245   : cube_lut_5 = 14'b10110011000110;
9'd246   : cube_lut_5 = 14'b10110011000111;
9'd247   : cube_lut_5 = 14'b10110011001000;
9'd248   : cube_lut_5 = 14'b10110011001010;
9'd249   : cube_lut_5 = 14'b10110011001011;
9'd250   : cube_lut_5 = 14'b10110011001100;
9'd251   : cube_lut_5 = 14'b10110011001110;
9'd252   : cube_lut_5 = 14'b10110011001111;
9'd253   : cube_lut_5 = 14'b10110011010001;
9'd254   : cube_lut_5 = 14'b10110011010010;
9'd255   : cube_lut_5 = 14'b10110011010011;
9'd256   : cube_lut_5 = 14'b10110011010101;
9'd257   : cube_lut_5 = 14'b10110011010110;
9'd258   : cube_lut_5 = 14'b10110011010111;
9'd259   : cube_lut_5 = 14'b10110011011001;
9'd260   : cube_lut_5 = 14'b10110011011010;
9'd261   : cube_lut_5 = 14'b10110011011011;
9'd262   : cube_lut_5 = 14'b10110011011101;
9'd263   : cube_lut_5 = 14'b10110011011110;
9'd264   : cube_lut_5 = 14'b10110011100000;
9'd265   : cube_lut_5 = 14'b10110011100001;
9'd266   : cube_lut_5 = 14'b10110011100010;
9'd267   : cube_lut_5 = 14'b10110011100100;
9'd268   : cube_lut_5 = 14'b10110011100101;
9'd269   : cube_lut_5 = 14'b10110011100110;
9'd270   : cube_lut_5 = 14'b10110011101000;
9'd271   : cube_lut_5 = 14'b10110011101001;
9'd272   : cube_lut_5 = 14'b10110011101010;
9'd273   : cube_lut_5 = 14'b10110011101100;
9'd274   : cube_lut_5 = 14'b10110011101101;
9'd275   : cube_lut_5 = 14'b10110011101110;
9'd276   : cube_lut_5 = 14'b10110011110000;
9'd277   : cube_lut_5 = 14'b10110011110001;
9'd278   : cube_lut_5 = 14'b10110011110010;
9'd279   : cube_lut_5 = 14'b10110011110100;
9'd280   : cube_lut_5 = 14'b10110011110101;
9'd281   : cube_lut_5 = 14'b10110011110111;
9'd282   : cube_lut_5 = 14'b10110011111000;
9'd283   : cube_lut_5 = 14'b10110011111001;
9'd284   : cube_lut_5 = 14'b10110011111011;
9'd285   : cube_lut_5 = 14'b10110011111100;
9'd286   : cube_lut_5 = 14'b10110011111101;
9'd287   : cube_lut_5 = 14'b10110011111111;
9'd288   : cube_lut_5 = 14'b10110100000000;
9'd289   : cube_lut_5 = 14'b10110100000001;
9'd290   : cube_lut_5 = 14'b10110100000011;
9'd291   : cube_lut_5 = 14'b10110100000100;
9'd292   : cube_lut_5 = 14'b10110100000101;
9'd293   : cube_lut_5 = 14'b10110100000111;
9'd294   : cube_lut_5 = 14'b10110100001000;
9'd295   : cube_lut_5 = 14'b10110100001001;
9'd296   : cube_lut_5 = 14'b10110100001011;
9'd297   : cube_lut_5 = 14'b10110100001100;
9'd298   : cube_lut_5 = 14'b10110100001101;
9'd299   : cube_lut_5 = 14'b10110100001111;
9'd300   : cube_lut_5 = 14'b10110100010000;
9'd301   : cube_lut_5 = 14'b10110100010001;
9'd302   : cube_lut_5 = 14'b10110100010011;
9'd303   : cube_lut_5 = 14'b10110100010100;
9'd304   : cube_lut_5 = 14'b10110100010101;
9'd305   : cube_lut_5 = 14'b10110100010111;
9'd306   : cube_lut_5 = 14'b10110100011000;
9'd307   : cube_lut_5 = 14'b10110100011010;
9'd308   : cube_lut_5 = 14'b10110100011011;
9'd309   : cube_lut_5 = 14'b10110100011100;
9'd310   : cube_lut_5 = 14'b10110100011110;
9'd311   : cube_lut_5 = 14'b10110100011111;
9'd312   : cube_lut_5 = 14'b10110100100000;
9'd313   : cube_lut_5 = 14'b10110100100010;
9'd314   : cube_lut_5 = 14'b10110100100011;
9'd315   : cube_lut_5 = 14'b10110100100100;
9'd316   : cube_lut_5 = 14'b10110100100110;
9'd317   : cube_lut_5 = 14'b10110100100111;
9'd318   : cube_lut_5 = 14'b10110100101000;
9'd319   : cube_lut_5 = 14'b10110100101010;
9'd320   : cube_lut_5 = 14'b10110100101011;
9'd321   : cube_lut_5 = 14'b10110100101100;
9'd322   : cube_lut_5 = 14'b10110100101110;
9'd323   : cube_lut_5 = 14'b10110100101111;
9'd324   : cube_lut_5 = 14'b10110100110000;
9'd325   : cube_lut_5 = 14'b10110100110010;
9'd326   : cube_lut_5 = 14'b10110100110011;
9'd327   : cube_lut_5 = 14'b10110100110100;
9'd328   : cube_lut_5 = 14'b10110100110110;
9'd329   : cube_lut_5 = 14'b10110100110111;
9'd330   : cube_lut_5 = 14'b10110100111000;
9'd331   : cube_lut_5 = 14'b10110100111010;
9'd332   : cube_lut_5 = 14'b10110100111011;
9'd333   : cube_lut_5 = 14'b10110100111100;
9'd334   : cube_lut_5 = 14'b10110100111110;
9'd335   : cube_lut_5 = 14'b10110100111111;
9'd336   : cube_lut_5 = 14'b10110101000000;
9'd337   : cube_lut_5 = 14'b10110101000010;
9'd338   : cube_lut_5 = 14'b10110101000011;
9'd339   : cube_lut_5 = 14'b10110101000100;
9'd340   : cube_lut_5 = 14'b10110101000110;
9'd341   : cube_lut_5 = 14'b10110101000111;
9'd342   : cube_lut_5 = 14'b10110101001000;
9'd343   : cube_lut_5 = 14'b10110101001010;
9'd344   : cube_lut_5 = 14'b10110101001011;
9'd345   : cube_lut_5 = 14'b10110101001100;
9'd346   : cube_lut_5 = 14'b10110101001110;
9'd347   : cube_lut_5 = 14'b10110101001111;
9'd348   : cube_lut_5 = 14'b10110101010000;
9'd349   : cube_lut_5 = 14'b10110101010010;
9'd350   : cube_lut_5 = 14'b10110101010011;
9'd351   : cube_lut_5 = 14'b10110101010100;
9'd352   : cube_lut_5 = 14'b10110101010110;
9'd353   : cube_lut_5 = 14'b10110101010111;
9'd354   : cube_lut_5 = 14'b10110101011000;
9'd355   : cube_lut_5 = 14'b10110101011010;
9'd356   : cube_lut_5 = 14'b10110101011011;
9'd357   : cube_lut_5 = 14'b10110101011100;
9'd358   : cube_lut_5 = 14'b10110101011110;
9'd359   : cube_lut_5 = 14'b10110101011111;
9'd360   : cube_lut_5 = 14'b10110101100000;
9'd361   : cube_lut_5 = 14'b10110101100010;
9'd362   : cube_lut_5 = 14'b10110101100011;
9'd363   : cube_lut_5 = 14'b10110101100100;
9'd364   : cube_lut_5 = 14'b10110101100110;
9'd365   : cube_lut_5 = 14'b10110101100111;
9'd366   : cube_lut_5 = 14'b10110101101000;
9'd367   : cube_lut_5 = 14'b10110101101010;
9'd368   : cube_lut_5 = 14'b10110101101011;
9'd369   : cube_lut_5 = 14'b10110101101100;
9'd370   : cube_lut_5 = 14'b10110101101101;
9'd371   : cube_lut_5 = 14'b10110101101111;
9'd372   : cube_lut_5 = 14'b10110101110000;
9'd373   : cube_lut_5 = 14'b10110101110001;
9'd374   : cube_lut_5 = 14'b10110101110011;
9'd375   : cube_lut_5 = 14'b10110101110100;
9'd376   : cube_lut_5 = 14'b10110101110101;
9'd377   : cube_lut_5 = 14'b10110101110111;
9'd378   : cube_lut_5 = 14'b10110101111000;
9'd379   : cube_lut_5 = 14'b10110101111001;
9'd380   : cube_lut_5 = 14'b10110101111011;
9'd381   : cube_lut_5 = 14'b10110101111100;
9'd382   : cube_lut_5 = 14'b10110101111101;
9'd383   : cube_lut_5 = 14'b10110101111111;
9'd384   : cube_lut_5 = 14'b10110110000000;
9'd385   : cube_lut_5 = 14'b10110110000001;
9'd386   : cube_lut_5 = 14'b10110110000011;
9'd387   : cube_lut_5 = 14'b10110110000100;
9'd388   : cube_lut_5 = 14'b10110110000101;
9'd389   : cube_lut_5 = 14'b10110110000111;
9'd390   : cube_lut_5 = 14'b10110110001000;
9'd391   : cube_lut_5 = 14'b10110110001001;
9'd392   : cube_lut_5 = 14'b10110110001011;
9'd393   : cube_lut_5 = 14'b10110110001100;
9'd394   : cube_lut_5 = 14'b10110110001101;
9'd395   : cube_lut_5 = 14'b10110110001110;
9'd396   : cube_lut_5 = 14'b10110110010000;
9'd397   : cube_lut_5 = 14'b10110110010001;
9'd398   : cube_lut_5 = 14'b10110110010010;
9'd399   : cube_lut_5 = 14'b10110110010100;
9'd400   : cube_lut_5 = 14'b10110110010101;
9'd401   : cube_lut_5 = 14'b10110110010110;
9'd402   : cube_lut_5 = 14'b10110110011000;
9'd403   : cube_lut_5 = 14'b10110110011001;
9'd404   : cube_lut_5 = 14'b10110110011010;
9'd405   : cube_lut_5 = 14'b10110110011100;
9'd406   : cube_lut_5 = 14'b10110110011101;
9'd407   : cube_lut_5 = 14'b10110110011110;
9'd408   : cube_lut_5 = 14'b10110110100000;
9'd409   : cube_lut_5 = 14'b10110110100001;
9'd410   : cube_lut_5 = 14'b10110110100010;
9'd411   : cube_lut_5 = 14'b10110110100011;
9'd412   : cube_lut_5 = 14'b10110110100101;
9'd413   : cube_lut_5 = 14'b10110110100110;
9'd414   : cube_lut_5 = 14'b10110110100111;
9'd415   : cube_lut_5 = 14'b10110110101001;
9'd416   : cube_lut_5 = 14'b10110110101010;
9'd417   : cube_lut_5 = 14'b10110110101011;
9'd418   : cube_lut_5 = 14'b10110110101101;
9'd419   : cube_lut_5 = 14'b10110110101110;
9'd420   : cube_lut_5 = 14'b10110110101111;
9'd421   : cube_lut_5 = 14'b10110110110001;
9'd422   : cube_lut_5 = 14'b10110110110010;
9'd423   : cube_lut_5 = 14'b10110110110011;
9'd424   : cube_lut_5 = 14'b10110110110100;
9'd425   : cube_lut_5 = 14'b10110110110110;
9'd426   : cube_lut_5 = 14'b10110110110111;
9'd427   : cube_lut_5 = 14'b10110110111000;
9'd428   : cube_lut_5 = 14'b10110110111010;
9'd429   : cube_lut_5 = 14'b10110110111011;
9'd430   : cube_lut_5 = 14'b10110110111100;
9'd431   : cube_lut_5 = 14'b10110110111110;
9'd432   : cube_lut_5 = 14'b10110110111111;
9'd433   : cube_lut_5 = 14'b10110111000000;
9'd434   : cube_lut_5 = 14'b10110111000010;
9'd435   : cube_lut_5 = 14'b10110111000011;
9'd436   : cube_lut_5 = 14'b10110111000100;
9'd437   : cube_lut_5 = 14'b10110111000101;
9'd438   : cube_lut_5 = 14'b10110111000111;
9'd439   : cube_lut_5 = 14'b10110111001000;
9'd440   : cube_lut_5 = 14'b10110111001001;
9'd441   : cube_lut_5 = 14'b10110111001011;
9'd442   : cube_lut_5 = 14'b10110111001100;
9'd443   : cube_lut_5 = 14'b10110111001101;
9'd444   : cube_lut_5 = 14'b10110111001111;
9'd445   : cube_lut_5 = 14'b10110111010000;
9'd446   : cube_lut_5 = 14'b10110111010001;
9'd447   : cube_lut_5 = 14'b10110111010010;
9'd448   : cube_lut_5 = 14'b10110111010100;
9'd449   : cube_lut_5 = 14'b10110111010101;
9'd450   : cube_lut_5 = 14'b10110111010110;
9'd451   : cube_lut_5 = 14'b10110111011000;
9'd452   : cube_lut_5 = 14'b10110111011001;
9'd453   : cube_lut_5 = 14'b10110111011010;
9'd454   : cube_lut_5 = 14'b10110111011100;
9'd455   : cube_lut_5 = 14'b10110111011101;
9'd456   : cube_lut_5 = 14'b10110111011110;
9'd457   : cube_lut_5 = 14'b10110111011111;
9'd458   : cube_lut_5 = 14'b10110111100001;
9'd459   : cube_lut_5 = 14'b10110111100010;
9'd460   : cube_lut_5 = 14'b10110111100011;
9'd461   : cube_lut_5 = 14'b10110111100101;
9'd462   : cube_lut_5 = 14'b10110111100110;
9'd463   : cube_lut_5 = 14'b10110111100111;
9'd464   : cube_lut_5 = 14'b10110111101001;
9'd465   : cube_lut_5 = 14'b10110111101010;
9'd466   : cube_lut_5 = 14'b10110111101011;
9'd467   : cube_lut_5 = 14'b10110111101100;
9'd468   : cube_lut_5 = 14'b10110111101110;
9'd469   : cube_lut_5 = 14'b10110111101111;
9'd470   : cube_lut_5 = 14'b10110111110000;
9'd471   : cube_lut_5 = 14'b10110111110010;
9'd472   : cube_lut_5 = 14'b10110111110011;
9'd473   : cube_lut_5 = 14'b10110111110100;
9'd474   : cube_lut_5 = 14'b10110111110101;
9'd475   : cube_lut_5 = 14'b10110111110111;
9'd476   : cube_lut_5 = 14'b10110111111000;
9'd477   : cube_lut_5 = 14'b10110111111001;
9'd478   : cube_lut_5 = 14'b10110111111011;
9'd479   : cube_lut_5 = 14'b10110111111100;
9'd480   : cube_lut_5 = 14'b10110111111101;
9'd481   : cube_lut_5 = 14'b10110111111111;
9'd482   : cube_lut_5 = 14'b10111000000000;
9'd483   : cube_lut_5 = 14'b10111000000001;
9'd484   : cube_lut_5 = 14'b10111000000010;
9'd485   : cube_lut_5 = 14'b10111000000100;
9'd486   : cube_lut_5 = 14'b10111000000101;
9'd487   : cube_lut_5 = 14'b10111000000110;
9'd488   : cube_lut_5 = 14'b10111000001000;
9'd489   : cube_lut_5 = 14'b10111000001001;
9'd490   : cube_lut_5 = 14'b10111000001010;
9'd491   : cube_lut_5 = 14'b10111000001011;
9'd492   : cube_lut_5 = 14'b10111000001101;
9'd493   : cube_lut_5 = 14'b10111000001110;
9'd494   : cube_lut_5 = 14'b10111000001111;
9'd495   : cube_lut_5 = 14'b10111000010001;
9'd496   : cube_lut_5 = 14'b10111000010010;
9'd497   : cube_lut_5 = 14'b10111000010011;
9'd498   : cube_lut_5 = 14'b10111000010100;
9'd499   : cube_lut_5 = 14'b10111000010110;
9'd500   : cube_lut_5 = 14'b10111000010111;
9'd501   : cube_lut_5 = 14'b10111000011000;
9'd502   : cube_lut_5 = 14'b10111000011010;
9'd503   : cube_lut_5 = 14'b10111000011011;
9'd504   : cube_lut_5 = 14'b10111000011100;
9'd505   : cube_lut_5 = 14'b10111000011101;
9'd506   : cube_lut_5 = 14'b10111000011111;
9'd507   : cube_lut_5 = 14'b10111000100000;
9'd508   : cube_lut_5 = 14'b10111000100001;
9'd509   : cube_lut_5 = 14'b10111000100011;
9'd510   : cube_lut_5 = 14'b10111000100100;
9'd511   : cube_lut_5 = 14'b10111000100101;

    endcase
end

always@* begin
    
    cube_lut_6 = 0;
    
    case(i_data[8:0])
 
 9'd0   : cube_lut_6 = 14'b10111000100110;
9'd1   : cube_lut_6 = 14'b10111000101000;
9'd2   : cube_lut_6 = 14'b10111000101001;
9'd3   : cube_lut_6 = 14'b10111000101010;
9'd4   : cube_lut_6 = 14'b10111000101100;
9'd5   : cube_lut_6 = 14'b10111000101101;
9'd6   : cube_lut_6 = 14'b10111000101110;
9'd7   : cube_lut_6 = 14'b10111000101111;
9'd8   : cube_lut_6 = 14'b10111000110001;
9'd9   : cube_lut_6 = 14'b10111000110010;
9'd10   : cube_lut_6 = 14'b10111000110011;
9'd11   : cube_lut_6 = 14'b10111000110100;
9'd12   : cube_lut_6 = 14'b10111000110110;
9'd13   : cube_lut_6 = 14'b10111000110111;
9'd14   : cube_lut_6 = 14'b10111000111000;
9'd15   : cube_lut_6 = 14'b10111000111010;
9'd16   : cube_lut_6 = 14'b10111000111011;
9'd17   : cube_lut_6 = 14'b10111000111100;
9'd18   : cube_lut_6 = 14'b10111000111101;
9'd19   : cube_lut_6 = 14'b10111000111111;
9'd20   : cube_lut_6 = 14'b10111001000000;
9'd21   : cube_lut_6 = 14'b10111001000001;
9'd22   : cube_lut_6 = 14'b10111001000011;
9'd23   : cube_lut_6 = 14'b10111001000100;
9'd24   : cube_lut_6 = 14'b10111001000101;
9'd25   : cube_lut_6 = 14'b10111001000110;
9'd26   : cube_lut_6 = 14'b10111001001000;
9'd27   : cube_lut_6 = 14'b10111001001001;
9'd28   : cube_lut_6 = 14'b10111001001010;
9'd29   : cube_lut_6 = 14'b10111001001011;
9'd30   : cube_lut_6 = 14'b10111001001101;
9'd31   : cube_lut_6 = 14'b10111001001110;
9'd32   : cube_lut_6 = 14'b10111001001111;
9'd33   : cube_lut_6 = 14'b10111001010001;
9'd34   : cube_lut_6 = 14'b10111001010010;
9'd35   : cube_lut_6 = 14'b10111001010011;
9'd36   : cube_lut_6 = 14'b10111001010100;
9'd37   : cube_lut_6 = 14'b10111001010110;
9'd38   : cube_lut_6 = 14'b10111001010111;
9'd39   : cube_lut_6 = 14'b10111001011000;
9'd40   : cube_lut_6 = 14'b10111001011001;
9'd41   : cube_lut_6 = 14'b10111001011011;
9'd42   : cube_lut_6 = 14'b10111001011100;
9'd43   : cube_lut_6 = 14'b10111001011101;
9'd44   : cube_lut_6 = 14'b10111001011111;
9'd45   : cube_lut_6 = 14'b10111001100000;
9'd46   : cube_lut_6 = 14'b10111001100001;
9'd47   : cube_lut_6 = 14'b10111001100010;
9'd48   : cube_lut_6 = 14'b10111001100100;
9'd49   : cube_lut_6 = 14'b10111001100101;
9'd50   : cube_lut_6 = 14'b10111001100110;
9'd51   : cube_lut_6 = 14'b10111001100111;
9'd52   : cube_lut_6 = 14'b10111001101001;
9'd53   : cube_lut_6 = 14'b10111001101010;
9'd54   : cube_lut_6 = 14'b10111001101011;
9'd55   : cube_lut_6 = 14'b10111001101101;
9'd56   : cube_lut_6 = 14'b10111001101110;
9'd57   : cube_lut_6 = 14'b10111001101111;
9'd58   : cube_lut_6 = 14'b10111001110000;
9'd59   : cube_lut_6 = 14'b10111001110010;
9'd60   : cube_lut_6 = 14'b10111001110011;
9'd61   : cube_lut_6 = 14'b10111001110100;
9'd62   : cube_lut_6 = 14'b10111001110101;
9'd63   : cube_lut_6 = 14'b10111001110111;
9'd64   : cube_lut_6 = 14'b10111001111000;
9'd65   : cube_lut_6 = 14'b10111001111001;
9'd66   : cube_lut_6 = 14'b10111001111010;
9'd67   : cube_lut_6 = 14'b10111001111100;
9'd68   : cube_lut_6 = 14'b10111001111101;
9'd69   : cube_lut_6 = 14'b10111001111110;
9'd70   : cube_lut_6 = 14'b10111001111111;
9'd71   : cube_lut_6 = 14'b10111010000001;
9'd72   : cube_lut_6 = 14'b10111010000010;
9'd73   : cube_lut_6 = 14'b10111010000011;
9'd74   : cube_lut_6 = 14'b10111010000101;
9'd75   : cube_lut_6 = 14'b10111010000110;
9'd76   : cube_lut_6 = 14'b10111010000111;
9'd77   : cube_lut_6 = 14'b10111010001000;
9'd78   : cube_lut_6 = 14'b10111010001010;
9'd79   : cube_lut_6 = 14'b10111010001011;
9'd80   : cube_lut_6 = 14'b10111010001100;
9'd81   : cube_lut_6 = 14'b10111010001101;
9'd82   : cube_lut_6 = 14'b10111010001111;
9'd83   : cube_lut_6 = 14'b10111010010000;
9'd84   : cube_lut_6 = 14'b10111010010001;
9'd85   : cube_lut_6 = 14'b10111010010010;
9'd86   : cube_lut_6 = 14'b10111010010100;
9'd87   : cube_lut_6 = 14'b10111010010101;
9'd88   : cube_lut_6 = 14'b10111010010110;
9'd89   : cube_lut_6 = 14'b10111010010111;
9'd90   : cube_lut_6 = 14'b10111010011001;
9'd91   : cube_lut_6 = 14'b10111010011010;
9'd92   : cube_lut_6 = 14'b10111010011011;
9'd93   : cube_lut_6 = 14'b10111010011100;
9'd94   : cube_lut_6 = 14'b10111010011110;
9'd95   : cube_lut_6 = 14'b10111010011111;
9'd96   : cube_lut_6 = 14'b10111010100000;
9'd97   : cube_lut_6 = 14'b10111010100001;
9'd98   : cube_lut_6 = 14'b10111010100011;
9'd99   : cube_lut_6 = 14'b10111010100100;
9'd100   : cube_lut_6 = 14'b10111010100101;
9'd101   : cube_lut_6 = 14'b10111010100110;
9'd102   : cube_lut_6 = 14'b10111010101000;
9'd103   : cube_lut_6 = 14'b10111010101001;
9'd104   : cube_lut_6 = 14'b10111010101010;
9'd105   : cube_lut_6 = 14'b10111010101100;
9'd106   : cube_lut_6 = 14'b10111010101101;
9'd107   : cube_lut_6 = 14'b10111010101110;
9'd108   : cube_lut_6 = 14'b10111010101111;
9'd109   : cube_lut_6 = 14'b10111010110001;
9'd110   : cube_lut_6 = 14'b10111010110010;
9'd111   : cube_lut_6 = 14'b10111010110011;
9'd112   : cube_lut_6 = 14'b10111010110100;
9'd113   : cube_lut_6 = 14'b10111010110110;
9'd114   : cube_lut_6 = 14'b10111010110111;
9'd115   : cube_lut_6 = 14'b10111010111000;
9'd116   : cube_lut_6 = 14'b10111010111001;
9'd117   : cube_lut_6 = 14'b10111010111011;
9'd118   : cube_lut_6 = 14'b10111010111100;
9'd119   : cube_lut_6 = 14'b10111010111101;
9'd120   : cube_lut_6 = 14'b10111010111110;
9'd121   : cube_lut_6 = 14'b10111011000000;
9'd122   : cube_lut_6 = 14'b10111011000001;
9'd123   : cube_lut_6 = 14'b10111011000010;
9'd124   : cube_lut_6 = 14'b10111011000011;
9'd125   : cube_lut_6 = 14'b10111011000101;
9'd126   : cube_lut_6 = 14'b10111011000110;
9'd127   : cube_lut_6 = 14'b10111011000111;
9'd128   : cube_lut_6 = 14'b10111011001000;
9'd129   : cube_lut_6 = 14'b10111011001010;
9'd130   : cube_lut_6 = 14'b10111011001011;
9'd131   : cube_lut_6 = 14'b10111011001100;
9'd132   : cube_lut_6 = 14'b10111011001101;
9'd133   : cube_lut_6 = 14'b10111011001111;
9'd134   : cube_lut_6 = 14'b10111011010000;
9'd135   : cube_lut_6 = 14'b10111011010001;
9'd136   : cube_lut_6 = 14'b10111011010010;
9'd137   : cube_lut_6 = 14'b10111011010011;
9'd138   : cube_lut_6 = 14'b10111011010101;
9'd139   : cube_lut_6 = 14'b10111011010110;
9'd140   : cube_lut_6 = 14'b10111011010111;
9'd141   : cube_lut_6 = 14'b10111011011000;
9'd142   : cube_lut_6 = 14'b10111011011010;
9'd143   : cube_lut_6 = 14'b10111011011011;
9'd144   : cube_lut_6 = 14'b10111011011100;
9'd145   : cube_lut_6 = 14'b10111011011101;
9'd146   : cube_lut_6 = 14'b10111011011111;
9'd147   : cube_lut_6 = 14'b10111011100000;
9'd148   : cube_lut_6 = 14'b10111011100001;
9'd149   : cube_lut_6 = 14'b10111011100010;
9'd150   : cube_lut_6 = 14'b10111011100100;
9'd151   : cube_lut_6 = 14'b10111011100101;
9'd152   : cube_lut_6 = 14'b10111011100110;
9'd153   : cube_lut_6 = 14'b10111011100111;
9'd154   : cube_lut_6 = 14'b10111011101001;
9'd155   : cube_lut_6 = 14'b10111011101010;
9'd156   : cube_lut_6 = 14'b10111011101011;
9'd157   : cube_lut_6 = 14'b10111011101100;
9'd158   : cube_lut_6 = 14'b10111011101110;
9'd159   : cube_lut_6 = 14'b10111011101111;
9'd160   : cube_lut_6 = 14'b10111011110000;
9'd161   : cube_lut_6 = 14'b10111011110001;
9'd162   : cube_lut_6 = 14'b10111011110011;
9'd163   : cube_lut_6 = 14'b10111011110100;
9'd164   : cube_lut_6 = 14'b10111011110101;
9'd165   : cube_lut_6 = 14'b10111011110110;
9'd166   : cube_lut_6 = 14'b10111011110111;
9'd167   : cube_lut_6 = 14'b10111011111001;
9'd168   : cube_lut_6 = 14'b10111011111010;
9'd169   : cube_lut_6 = 14'b10111011111011;
9'd170   : cube_lut_6 = 14'b10111011111100;
9'd171   : cube_lut_6 = 14'b10111011111110;
9'd172   : cube_lut_6 = 14'b10111011111111;
9'd173   : cube_lut_6 = 14'b10111100000000;
9'd174   : cube_lut_6 = 14'b10111100000001;
9'd175   : cube_lut_6 = 14'b10111100000011;
9'd176   : cube_lut_6 = 14'b10111100000100;
9'd177   : cube_lut_6 = 14'b10111100000101;
9'd178   : cube_lut_6 = 14'b10111100000110;
9'd179   : cube_lut_6 = 14'b10111100001000;
9'd180   : cube_lut_6 = 14'b10111100001001;
9'd181   : cube_lut_6 = 14'b10111100001010;
9'd182   : cube_lut_6 = 14'b10111100001011;
9'd183   : cube_lut_6 = 14'b10111100001101;
9'd184   : cube_lut_6 = 14'b10111100001110;
9'd185   : cube_lut_6 = 14'b10111100001111;
9'd186   : cube_lut_6 = 14'b10111100010000;
9'd187   : cube_lut_6 = 14'b10111100010001;
9'd188   : cube_lut_6 = 14'b10111100010011;
9'd189   : cube_lut_6 = 14'b10111100010100;
9'd190   : cube_lut_6 = 14'b10111100010101;
9'd191   : cube_lut_6 = 14'b10111100010110;
9'd192   : cube_lut_6 = 14'b10111100011000;
9'd193   : cube_lut_6 = 14'b10111100011001;
9'd194   : cube_lut_6 = 14'b10111100011010;
9'd195   : cube_lut_6 = 14'b10111100011011;
9'd196   : cube_lut_6 = 14'b10111100011101;
9'd197   : cube_lut_6 = 14'b10111100011110;
9'd198   : cube_lut_6 = 14'b10111100011111;
9'd199   : cube_lut_6 = 14'b10111100100000;
9'd200   : cube_lut_6 = 14'b10111100100001;
9'd201   : cube_lut_6 = 14'b10111100100011;
9'd202   : cube_lut_6 = 14'b10111100100100;
9'd203   : cube_lut_6 = 14'b10111100100101;
9'd204   : cube_lut_6 = 14'b10111100100110;
9'd205   : cube_lut_6 = 14'b10111100101000;
9'd206   : cube_lut_6 = 14'b10111100101001;
9'd207   : cube_lut_6 = 14'b10111100101010;
9'd208   : cube_lut_6 = 14'b10111100101011;
9'd209   : cube_lut_6 = 14'b10111100101100;
9'd210   : cube_lut_6 = 14'b10111100101110;
9'd211   : cube_lut_6 = 14'b10111100101111;
9'd212   : cube_lut_6 = 14'b10111100110000;
9'd213   : cube_lut_6 = 14'b10111100110001;
9'd214   : cube_lut_6 = 14'b10111100110011;
9'd215   : cube_lut_6 = 14'b10111100110100;
9'd216   : cube_lut_6 = 14'b10111100110101;
9'd217   : cube_lut_6 = 14'b10111100110110;
9'd218   : cube_lut_6 = 14'b10111100111000;
9'd219   : cube_lut_6 = 14'b10111100111001;
9'd220   : cube_lut_6 = 14'b10111100111010;
9'd221   : cube_lut_6 = 14'b10111100111011;
9'd222   : cube_lut_6 = 14'b10111100111100;
9'd223   : cube_lut_6 = 14'b10111100111110;
9'd224   : cube_lut_6 = 14'b10111100111111;
9'd225   : cube_lut_6 = 14'b10111101000000;
9'd226   : cube_lut_6 = 14'b10111101000001;
9'd227   : cube_lut_6 = 14'b10111101000011;
9'd228   : cube_lut_6 = 14'b10111101000100;
9'd229   : cube_lut_6 = 14'b10111101000101;
9'd230   : cube_lut_6 = 14'b10111101000110;
9'd231   : cube_lut_6 = 14'b10111101000111;
9'd232   : cube_lut_6 = 14'b10111101001001;
9'd233   : cube_lut_6 = 14'b10111101001010;
9'd234   : cube_lut_6 = 14'b10111101001011;
9'd235   : cube_lut_6 = 14'b10111101001100;
9'd236   : cube_lut_6 = 14'b10111101001110;
9'd237   : cube_lut_6 = 14'b10111101001111;
9'd238   : cube_lut_6 = 14'b10111101010000;
9'd239   : cube_lut_6 = 14'b10111101010001;
9'd240   : cube_lut_6 = 14'b10111101010010;
9'd241   : cube_lut_6 = 14'b10111101010100;
9'd242   : cube_lut_6 = 14'b10111101010101;
9'd243   : cube_lut_6 = 14'b10111101010110;
9'd244   : cube_lut_6 = 14'b10111101010111;
9'd245   : cube_lut_6 = 14'b10111101011000;
9'd246   : cube_lut_6 = 14'b10111101011010;
9'd247   : cube_lut_6 = 14'b10111101011011;
9'd248   : cube_lut_6 = 14'b10111101011100;
9'd249   : cube_lut_6 = 14'b10111101011101;
9'd250   : cube_lut_6 = 14'b10111101011111;
9'd251   : cube_lut_6 = 14'b10111101100000;
9'd252   : cube_lut_6 = 14'b10111101100001;
9'd253   : cube_lut_6 = 14'b10111101100010;
9'd254   : cube_lut_6 = 14'b10111101100011;
9'd255   : cube_lut_6 = 14'b10111101100101;
9'd256   : cube_lut_6 = 14'b10111101100110;
9'd257   : cube_lut_6 = 14'b10111101100111;
9'd258   : cube_lut_6 = 14'b10111101101000;
9'd259   : cube_lut_6 = 14'b10111101101010;
9'd260   : cube_lut_6 = 14'b10111101101011;
9'd261   : cube_lut_6 = 14'b10111101101100;
9'd262   : cube_lut_6 = 14'b10111101101101;
9'd263   : cube_lut_6 = 14'b10111101101110;
9'd264   : cube_lut_6 = 14'b10111101110000;
9'd265   : cube_lut_6 = 14'b10111101110001;
9'd266   : cube_lut_6 = 14'b10111101110010;
9'd267   : cube_lut_6 = 14'b10111101110011;
9'd268   : cube_lut_6 = 14'b10111101110100;
9'd269   : cube_lut_6 = 14'b10111101110110;
9'd270   : cube_lut_6 = 14'b10111101110111;
9'd271   : cube_lut_6 = 14'b10111101111000;
9'd272   : cube_lut_6 = 14'b10111101111001;
9'd273   : cube_lut_6 = 14'b10111101111011;
9'd274   : cube_lut_6 = 14'b10111101111100;
9'd275   : cube_lut_6 = 14'b10111101111101;
9'd276   : cube_lut_6 = 14'b10111101111110;
9'd277   : cube_lut_6 = 14'b10111101111111;
9'd278   : cube_lut_6 = 14'b10111110000001;
9'd279   : cube_lut_6 = 14'b10111110000010;
9'd280   : cube_lut_6 = 14'b10111110000011;
9'd281   : cube_lut_6 = 14'b10111110000100;
9'd282   : cube_lut_6 = 14'b10111110000101;
9'd283   : cube_lut_6 = 14'b10111110000111;
9'd284   : cube_lut_6 = 14'b10111110001000;
9'd285   : cube_lut_6 = 14'b10111110001001;
9'd286   : cube_lut_6 = 14'b10111110001010;
9'd287   : cube_lut_6 = 14'b10111110001011;
9'd288   : cube_lut_6 = 14'b10111110001101;
9'd289   : cube_lut_6 = 14'b10111110001110;
9'd290   : cube_lut_6 = 14'b10111110001111;
9'd291   : cube_lut_6 = 14'b10111110010000;
9'd292   : cube_lut_6 = 14'b10111110010001;
9'd293   : cube_lut_6 = 14'b10111110010011;
9'd294   : cube_lut_6 = 14'b10111110010100;
9'd295   : cube_lut_6 = 14'b10111110010101;
9'd296   : cube_lut_6 = 14'b10111110010110;
9'd297   : cube_lut_6 = 14'b10111110011000;
9'd298   : cube_lut_6 = 14'b10111110011001;
9'd299   : cube_lut_6 = 14'b10111110011010;
9'd300   : cube_lut_6 = 14'b10111110011011;
9'd301   : cube_lut_6 = 14'b10111110011100;
9'd302   : cube_lut_6 = 14'b10111110011110;
9'd303   : cube_lut_6 = 14'b10111110011111;
9'd304   : cube_lut_6 = 14'b10111110100000;
9'd305   : cube_lut_6 = 14'b10111110100001;
9'd306   : cube_lut_6 = 14'b10111110100010;
9'd307   : cube_lut_6 = 14'b10111110100100;
9'd308   : cube_lut_6 = 14'b10111110100101;
9'd309   : cube_lut_6 = 14'b10111110100110;
9'd310   : cube_lut_6 = 14'b10111110100111;
9'd311   : cube_lut_6 = 14'b10111110101000;
9'd312   : cube_lut_6 = 14'b10111110101010;
9'd313   : cube_lut_6 = 14'b10111110101011;
9'd314   : cube_lut_6 = 14'b10111110101100;
9'd315   : cube_lut_6 = 14'b10111110101101;
9'd316   : cube_lut_6 = 14'b10111110101110;
9'd317   : cube_lut_6 = 14'b10111110110000;
9'd318   : cube_lut_6 = 14'b10111110110001;
9'd319   : cube_lut_6 = 14'b10111110110010;
9'd320   : cube_lut_6 = 14'b10111110110011;
9'd321   : cube_lut_6 = 14'b10111110110100;
9'd322   : cube_lut_6 = 14'b10111110110110;
9'd323   : cube_lut_6 = 14'b10111110110111;
9'd324   : cube_lut_6 = 14'b10111110111000;
9'd325   : cube_lut_6 = 14'b10111110111001;
9'd326   : cube_lut_6 = 14'b10111110111010;
9'd327   : cube_lut_6 = 14'b10111110111100;
9'd328   : cube_lut_6 = 14'b10111110111101;
9'd329   : cube_lut_6 = 14'b10111110111110;
9'd330   : cube_lut_6 = 14'b10111110111111;
9'd331   : cube_lut_6 = 14'b10111111000000;
9'd332   : cube_lut_6 = 14'b10111111000010;
9'd333   : cube_lut_6 = 14'b10111111000011;
9'd334   : cube_lut_6 = 14'b10111111000100;
9'd335   : cube_lut_6 = 14'b10111111000101;
9'd336   : cube_lut_6 = 14'b10111111000110;
9'd337   : cube_lut_6 = 14'b10111111001000;
9'd338   : cube_lut_6 = 14'b10111111001001;
9'd339   : cube_lut_6 = 14'b10111111001010;
9'd340   : cube_lut_6 = 14'b10111111001011;
9'd341   : cube_lut_6 = 14'b10111111001100;
9'd342   : cube_lut_6 = 14'b10111111001110;
9'd343   : cube_lut_6 = 14'b10111111001111;
9'd344   : cube_lut_6 = 14'b10111111010000;
9'd345   : cube_lut_6 = 14'b10111111010001;
9'd346   : cube_lut_6 = 14'b10111111010010;
9'd347   : cube_lut_6 = 14'b10111111010011;
9'd348   : cube_lut_6 = 14'b10111111010101;
9'd349   : cube_lut_6 = 14'b10111111010110;
9'd350   : cube_lut_6 = 14'b10111111010111;
9'd351   : cube_lut_6 = 14'b10111111011000;
9'd352   : cube_lut_6 = 14'b10111111011001;
9'd353   : cube_lut_6 = 14'b10111111011011;
9'd354   : cube_lut_6 = 14'b10111111011100;
9'd355   : cube_lut_6 = 14'b10111111011101;
9'd356   : cube_lut_6 = 14'b10111111011110;
9'd357   : cube_lut_6 = 14'b10111111011111;
9'd358   : cube_lut_6 = 14'b10111111100001;
9'd359   : cube_lut_6 = 14'b10111111100010;
9'd360   : cube_lut_6 = 14'b10111111100011;
9'd361   : cube_lut_6 = 14'b10111111100100;
9'd362   : cube_lut_6 = 14'b10111111100101;
9'd363   : cube_lut_6 = 14'b10111111100111;
9'd364   : cube_lut_6 = 14'b10111111101000;
9'd365   : cube_lut_6 = 14'b10111111101001;
9'd366   : cube_lut_6 = 14'b10111111101010;
9'd367   : cube_lut_6 = 14'b10111111101011;
9'd368   : cube_lut_6 = 14'b10111111101101;
9'd369   : cube_lut_6 = 14'b10111111101110;
9'd370   : cube_lut_6 = 14'b10111111101111;
9'd371   : cube_lut_6 = 14'b10111111110000;
9'd372   : cube_lut_6 = 14'b10111111110001;
9'd373   : cube_lut_6 = 14'b10111111110010;
9'd374   : cube_lut_6 = 14'b10111111110100;
9'd375   : cube_lut_6 = 14'b10111111110101;
9'd376   : cube_lut_6 = 14'b10111111110110;
9'd377   : cube_lut_6 = 14'b10111111110111;
9'd378   : cube_lut_6 = 14'b10111111111000;
9'd379   : cube_lut_6 = 14'b10111111111010;
9'd380   : cube_lut_6 = 14'b10111111111011;
9'd381   : cube_lut_6 = 14'b10111111111100;
9'd382   : cube_lut_6 = 14'b10111111111101;
9'd383   : cube_lut_6 = 14'b10111111111110;
9'd384   : cube_lut_6 = 14'b11000000000000;
9'd385   : cube_lut_6 = 14'b11000000000001;
9'd386   : cube_lut_6 = 14'b11000000000010;
9'd387   : cube_lut_6 = 14'b11000000000011;
9'd388   : cube_lut_6 = 14'b11000000000100;
9'd389   : cube_lut_6 = 14'b11000000000101;
9'd390   : cube_lut_6 = 14'b11000000000111;
9'd391   : cube_lut_6 = 14'b11000000001000;
9'd392   : cube_lut_6 = 14'b11000000001001;
9'd393   : cube_lut_6 = 14'b11000000001010;
9'd394   : cube_lut_6 = 14'b11000000001011;
9'd395   : cube_lut_6 = 14'b11000000001101;
9'd396   : cube_lut_6 = 14'b11000000001110;
9'd397   : cube_lut_6 = 14'b11000000001111;
9'd398   : cube_lut_6 = 14'b11000000010000;
9'd399   : cube_lut_6 = 14'b11000000010001;
9'd400   : cube_lut_6 = 14'b11000000010010;
9'd401   : cube_lut_6 = 14'b11000000010100;
9'd402   : cube_lut_6 = 14'b11000000010101;
9'd403   : cube_lut_6 = 14'b11000000010110;
9'd404   : cube_lut_6 = 14'b11000000010111;
9'd405   : cube_lut_6 = 14'b11000000011000;
9'd406   : cube_lut_6 = 14'b11000000011010;
9'd407   : cube_lut_6 = 14'b11000000011011;
9'd408   : cube_lut_6 = 14'b11000000011100;
9'd409   : cube_lut_6 = 14'b11000000011101;
9'd410   : cube_lut_6 = 14'b11000000011110;
9'd411   : cube_lut_6 = 14'b11000000011111;
9'd412   : cube_lut_6 = 14'b11000000100001;
9'd413   : cube_lut_6 = 14'b11000000100010;
9'd414   : cube_lut_6 = 14'b11000000100011;
9'd415   : cube_lut_6 = 14'b11000000100100;
9'd416   : cube_lut_6 = 14'b11000000100101;
9'd417   : cube_lut_6 = 14'b11000000100110;
9'd418   : cube_lut_6 = 14'b11000000101000;
9'd419   : cube_lut_6 = 14'b11000000101001;
9'd420   : cube_lut_6 = 14'b11000000101010;
9'd421   : cube_lut_6 = 14'b11000000101011;
9'd422   : cube_lut_6 = 14'b11000000101100;
9'd423   : cube_lut_6 = 14'b11000000101110;
9'd424   : cube_lut_6 = 14'b11000000101111;
9'd425   : cube_lut_6 = 14'b11000000110000;
9'd426   : cube_lut_6 = 14'b11000000110001;
9'd427   : cube_lut_6 = 14'b11000000110010;
9'd428   : cube_lut_6 = 14'b11000000110011;
9'd429   : cube_lut_6 = 14'b11000000110101;
9'd430   : cube_lut_6 = 14'b11000000110110;
9'd431   : cube_lut_6 = 14'b11000000110111;
9'd432   : cube_lut_6 = 14'b11000000111000;
9'd433   : cube_lut_6 = 14'b11000000111001;
9'd434   : cube_lut_6 = 14'b11000000111010;
9'd435   : cube_lut_6 = 14'b11000000111100;
9'd436   : cube_lut_6 = 14'b11000000111101;
9'd437   : cube_lut_6 = 14'b11000000111110;
9'd438   : cube_lut_6 = 14'b11000000111111;
9'd439   : cube_lut_6 = 14'b11000001000000;
9'd440   : cube_lut_6 = 14'b11000001000010;
9'd441   : cube_lut_6 = 14'b11000001000011;
9'd442   : cube_lut_6 = 14'b11000001000100;
9'd443   : cube_lut_6 = 14'b11000001000101;
9'd444   : cube_lut_6 = 14'b11000001000110;
9'd445   : cube_lut_6 = 14'b11000001000111;
9'd446   : cube_lut_6 = 14'b11000001001001;
9'd447   : cube_lut_6 = 14'b11000001001010;
9'd448   : cube_lut_6 = 14'b11000001001011;
9'd449   : cube_lut_6 = 14'b11000001001100;
9'd450   : cube_lut_6 = 14'b11000001001101;
9'd451   : cube_lut_6 = 14'b11000001001110;
9'd452   : cube_lut_6 = 14'b11000001010000;
9'd453   : cube_lut_6 = 14'b11000001010001;
9'd454   : cube_lut_6 = 14'b11000001010010;
9'd455   : cube_lut_6 = 14'b11000001010011;
9'd456   : cube_lut_6 = 14'b11000001010100;
9'd457   : cube_lut_6 = 14'b11000001010101;
9'd458   : cube_lut_6 = 14'b11000001010111;
9'd459   : cube_lut_6 = 14'b11000001011000;
9'd460   : cube_lut_6 = 14'b11000001011001;
9'd461   : cube_lut_6 = 14'b11000001011010;
9'd462   : cube_lut_6 = 14'b11000001011011;
9'd463   : cube_lut_6 = 14'b11000001011100;
9'd464   : cube_lut_6 = 14'b11000001011110;
9'd465   : cube_lut_6 = 14'b11000001011111;
9'd466   : cube_lut_6 = 14'b11000001100000;
9'd467   : cube_lut_6 = 14'b11000001100001;
9'd468   : cube_lut_6 = 14'b11000001100010;
9'd469   : cube_lut_6 = 14'b11000001100011;
9'd470   : cube_lut_6 = 14'b11000001100101;
9'd471   : cube_lut_6 = 14'b11000001100110;
9'd472   : cube_lut_6 = 14'b11000001100111;
9'd473   : cube_lut_6 = 14'b11000001101000;
9'd474   : cube_lut_6 = 14'b11000001101001;
9'd475   : cube_lut_6 = 14'b11000001101010;
9'd476   : cube_lut_6 = 14'b11000001101100;
9'd477   : cube_lut_6 = 14'b11000001101101;
9'd478   : cube_lut_6 = 14'b11000001101110;
9'd479   : cube_lut_6 = 14'b11000001101111;
9'd480   : cube_lut_6 = 14'b11000001110000;
9'd481   : cube_lut_6 = 14'b11000001110001;
9'd482   : cube_lut_6 = 14'b11000001110011;
9'd483   : cube_lut_6 = 14'b11000001110100;
9'd484   : cube_lut_6 = 14'b11000001110101;
9'd485   : cube_lut_6 = 14'b11000001110110;
9'd486   : cube_lut_6 = 14'b11000001110111;
9'd487   : cube_lut_6 = 14'b11000001111000;
9'd488   : cube_lut_6 = 14'b11000001111010;
9'd489   : cube_lut_6 = 14'b11000001111011;
9'd490   : cube_lut_6 = 14'b11000001111100;
9'd491   : cube_lut_6 = 14'b11000001111101;
9'd492   : cube_lut_6 = 14'b11000001111110;
9'd493   : cube_lut_6 = 14'b11000001111111;
9'd494   : cube_lut_6 = 14'b11000010000001;
9'd495   : cube_lut_6 = 14'b11000010000010;
9'd496   : cube_lut_6 = 14'b11000010000011;
9'd497   : cube_lut_6 = 14'b11000010000100;
9'd498   : cube_lut_6 = 14'b11000010000101;
9'd499   : cube_lut_6 = 14'b11000010000110;
9'd500   : cube_lut_6 = 14'b11000010000111;
9'd501   : cube_lut_6 = 14'b11000010001001;
9'd502   : cube_lut_6 = 14'b11000010001010;
9'd503   : cube_lut_6 = 14'b11000010001011;
9'd504   : cube_lut_6 = 14'b11000010001100;
9'd505   : cube_lut_6 = 14'b11000010001101;
9'd506   : cube_lut_6 = 14'b11000010001110;
9'd507   : cube_lut_6 = 14'b11000010010000;
9'd508   : cube_lut_6 = 14'b11000010010001;
9'd509   : cube_lut_6 = 14'b11000010010010;
9'd510   : cube_lut_6 = 14'b11000010010011;
9'd511   : cube_lut_6 = 14'b11000010010100;

    endcase
end

always@* begin
    
    cube_lut_7 = 0;
    
    case(i_data[8:0])
 
 9'd0   : cube_lut_7 = 14'b11000010010101;
9'd1   : cube_lut_7 = 14'b11000010010111;
9'd2   : cube_lut_7 = 14'b11000010011000;
9'd3   : cube_lut_7 = 14'b11000010011001;
9'd4   : cube_lut_7 = 14'b11000010011010;
9'd5   : cube_lut_7 = 14'b11000010011011;
9'd6   : cube_lut_7 = 14'b11000010011100;
9'd7   : cube_lut_7 = 14'b11000010011101;
9'd8   : cube_lut_7 = 14'b11000010011111;
9'd9   : cube_lut_7 = 14'b11000010100000;
9'd10   : cube_lut_7 = 14'b11000010100001;
9'd11   : cube_lut_7 = 14'b11000010100010;
9'd12   : cube_lut_7 = 14'b11000010100011;
9'd13   : cube_lut_7 = 14'b11000010100100;
9'd14   : cube_lut_7 = 14'b11000010100110;
9'd15   : cube_lut_7 = 14'b11000010100111;
9'd16   : cube_lut_7 = 14'b11000010101000;
9'd17   : cube_lut_7 = 14'b11000010101001;
9'd18   : cube_lut_7 = 14'b11000010101010;
9'd19   : cube_lut_7 = 14'b11000010101011;
9'd20   : cube_lut_7 = 14'b11000010101100;
9'd21   : cube_lut_7 = 14'b11000010101110;
9'd22   : cube_lut_7 = 14'b11000010101111;
9'd23   : cube_lut_7 = 14'b11000010110000;
9'd24   : cube_lut_7 = 14'b11000010110001;
9'd25   : cube_lut_7 = 14'b11000010110010;
9'd26   : cube_lut_7 = 14'b11000010110011;
9'd27   : cube_lut_7 = 14'b11000010110101;
9'd28   : cube_lut_7 = 14'b11000010110110;
9'd29   : cube_lut_7 = 14'b11000010110111;
9'd30   : cube_lut_7 = 14'b11000010111000;
9'd31   : cube_lut_7 = 14'b11000010111001;
9'd32   : cube_lut_7 = 14'b11000010111010;
9'd33   : cube_lut_7 = 14'b11000010111011;
9'd34   : cube_lut_7 = 14'b11000010111101;
9'd35   : cube_lut_7 = 14'b11000010111110;
9'd36   : cube_lut_7 = 14'b11000010111111;
9'd37   : cube_lut_7 = 14'b11000011000000;
9'd38   : cube_lut_7 = 14'b11000011000001;
9'd39   : cube_lut_7 = 14'b11000011000010;
9'd40   : cube_lut_7 = 14'b11000011000011;
9'd41   : cube_lut_7 = 14'b11000011000101;
9'd42   : cube_lut_7 = 14'b11000011000110;
9'd43   : cube_lut_7 = 14'b11000011000111;
9'd44   : cube_lut_7 = 14'b11000011001000;
9'd45   : cube_lut_7 = 14'b11000011001001;
9'd46   : cube_lut_7 = 14'b11000011001010;
9'd47   : cube_lut_7 = 14'b11000011001100;
9'd48   : cube_lut_7 = 14'b11000011001101;
9'd49   : cube_lut_7 = 14'b11000011001110;
9'd50   : cube_lut_7 = 14'b11000011001111;
9'd51   : cube_lut_7 = 14'b11000011010000;
9'd52   : cube_lut_7 = 14'b11000011010001;
9'd53   : cube_lut_7 = 14'b11000011010010;
9'd54   : cube_lut_7 = 14'b11000011010100;
9'd55   : cube_lut_7 = 14'b11000011010101;
9'd56   : cube_lut_7 = 14'b11000011010110;
9'd57   : cube_lut_7 = 14'b11000011010111;
9'd58   : cube_lut_7 = 14'b11000011011000;
9'd59   : cube_lut_7 = 14'b11000011011001;
9'd60   : cube_lut_7 = 14'b11000011011010;
9'd61   : cube_lut_7 = 14'b11000011011100;
9'd62   : cube_lut_7 = 14'b11000011011101;
9'd63   : cube_lut_7 = 14'b11000011011110;
9'd64   : cube_lut_7 = 14'b11000011011111;
9'd65   : cube_lut_7 = 14'b11000011100000;
9'd66   : cube_lut_7 = 14'b11000011100001;
9'd67   : cube_lut_7 = 14'b11000011100010;
9'd68   : cube_lut_7 = 14'b11000011100100;
9'd69   : cube_lut_7 = 14'b11000011100101;
9'd70   : cube_lut_7 = 14'b11000011100110;
9'd71   : cube_lut_7 = 14'b11000011100111;
9'd72   : cube_lut_7 = 14'b11000011101000;
9'd73   : cube_lut_7 = 14'b11000011101001;
9'd74   : cube_lut_7 = 14'b11000011101010;
9'd75   : cube_lut_7 = 14'b11000011101100;
9'd76   : cube_lut_7 = 14'b11000011101101;
9'd77   : cube_lut_7 = 14'b11000011101110;
9'd78   : cube_lut_7 = 14'b11000011101111;
9'd79   : cube_lut_7 = 14'b11000011110000;
9'd80   : cube_lut_7 = 14'b11000011110001;
9'd81   : cube_lut_7 = 14'b11000011110010;
9'd82   : cube_lut_7 = 14'b11000011110100;
9'd83   : cube_lut_7 = 14'b11000011110101;
9'd84   : cube_lut_7 = 14'b11000011110110;
9'd85   : cube_lut_7 = 14'b11000011110111;
9'd86   : cube_lut_7 = 14'b11000011111000;
9'd87   : cube_lut_7 = 14'b11000011111001;
9'd88   : cube_lut_7 = 14'b11000011111010;
9'd89   : cube_lut_7 = 14'b11000011111011;
9'd90   : cube_lut_7 = 14'b11000011111101;
9'd91   : cube_lut_7 = 14'b11000011111110;
9'd92   : cube_lut_7 = 14'b11000011111111;
9'd93   : cube_lut_7 = 14'b11000100000000;
9'd94   : cube_lut_7 = 14'b11000100000001;
9'd95   : cube_lut_7 = 14'b11000100000010;
9'd96   : cube_lut_7 = 14'b11000100000011;
9'd97   : cube_lut_7 = 14'b11000100000101;
9'd98   : cube_lut_7 = 14'b11000100000110;
9'd99   : cube_lut_7 = 14'b11000100000111;
9'd100   : cube_lut_7 = 14'b11000100001000;
9'd101   : cube_lut_7 = 14'b11000100001001;
9'd102   : cube_lut_7 = 14'b11000100001010;
9'd103   : cube_lut_7 = 14'b11000100001011;
9'd104   : cube_lut_7 = 14'b11000100001101;
9'd105   : cube_lut_7 = 14'b11000100001110;
9'd106   : cube_lut_7 = 14'b11000100001111;
9'd107   : cube_lut_7 = 14'b11000100010000;
9'd108   : cube_lut_7 = 14'b11000100010001;
9'd109   : cube_lut_7 = 14'b11000100010010;
9'd110   : cube_lut_7 = 14'b11000100010011;
9'd111   : cube_lut_7 = 14'b11000100010100;
9'd112   : cube_lut_7 = 14'b11000100010110;
9'd113   : cube_lut_7 = 14'b11000100010111;
9'd114   : cube_lut_7 = 14'b11000100011000;
9'd115   : cube_lut_7 = 14'b11000100011001;
9'd116   : cube_lut_7 = 14'b11000100011010;
9'd117   : cube_lut_7 = 14'b11000100011011;
9'd118   : cube_lut_7 = 14'b11000100011100;
9'd119   : cube_lut_7 = 14'b11000100011110;
9'd120   : cube_lut_7 = 14'b11000100011111;
9'd121   : cube_lut_7 = 14'b11000100100000;
9'd122   : cube_lut_7 = 14'b11000100100001;
9'd123   : cube_lut_7 = 14'b11000100100010;
9'd124   : cube_lut_7 = 14'b11000100100011;
9'd125   : cube_lut_7 = 14'b11000100100100;
9'd126   : cube_lut_7 = 14'b11000100100101;
9'd127   : cube_lut_7 = 14'b11000100100111;
9'd128   : cube_lut_7 = 14'b11000100101000;
9'd129   : cube_lut_7 = 14'b11000100101001;
9'd130   : cube_lut_7 = 14'b11000100101010;
9'd131   : cube_lut_7 = 14'b11000100101011;
9'd132   : cube_lut_7 = 14'b11000100101100;
9'd133   : cube_lut_7 = 14'b11000100101101;
9'd134   : cube_lut_7 = 14'b11000100101110;
9'd135   : cube_lut_7 = 14'b11000100110000;
9'd136   : cube_lut_7 = 14'b11000100110001;
9'd137   : cube_lut_7 = 14'b11000100110010;
9'd138   : cube_lut_7 = 14'b11000100110011;
9'd139   : cube_lut_7 = 14'b11000100110100;
9'd140   : cube_lut_7 = 14'b11000100110101;
9'd141   : cube_lut_7 = 14'b11000100110110;
9'd142   : cube_lut_7 = 14'b11000100111000;
9'd143   : cube_lut_7 = 14'b11000100111001;
9'd144   : cube_lut_7 = 14'b11000100111010;
9'd145   : cube_lut_7 = 14'b11000100111011;
9'd146   : cube_lut_7 = 14'b11000100111100;
9'd147   : cube_lut_7 = 14'b11000100111101;
9'd148   : cube_lut_7 = 14'b11000100111110;
9'd149   : cube_lut_7 = 14'b11000100111111;
9'd150   : cube_lut_7 = 14'b11000101000001;
9'd151   : cube_lut_7 = 14'b11000101000010;
9'd152   : cube_lut_7 = 14'b11000101000011;
9'd153   : cube_lut_7 = 14'b11000101000100;
9'd154   : cube_lut_7 = 14'b11000101000101;
9'd155   : cube_lut_7 = 14'b11000101000110;
9'd156   : cube_lut_7 = 14'b11000101000111;
9'd157   : cube_lut_7 = 14'b11000101001000;
9'd158   : cube_lut_7 = 14'b11000101001010;
9'd159   : cube_lut_7 = 14'b11000101001011;
9'd160   : cube_lut_7 = 14'b11000101001100;
9'd161   : cube_lut_7 = 14'b11000101001101;
9'd162   : cube_lut_7 = 14'b11000101001110;
9'd163   : cube_lut_7 = 14'b11000101001111;
9'd164   : cube_lut_7 = 14'b11000101010000;
9'd165   : cube_lut_7 = 14'b11000101010001;
9'd166   : cube_lut_7 = 14'b11000101010011;
9'd167   : cube_lut_7 = 14'b11000101010100;
9'd168   : cube_lut_7 = 14'b11000101010101;
9'd169   : cube_lut_7 = 14'b11000101010110;
9'd170   : cube_lut_7 = 14'b11000101010111;
9'd171   : cube_lut_7 = 14'b11000101011000;
9'd172   : cube_lut_7 = 14'b11000101011001;
9'd173   : cube_lut_7 = 14'b11000101011010;
9'd174   : cube_lut_7 = 14'b11000101011011;
9'd175   : cube_lut_7 = 14'b11000101011101;
9'd176   : cube_lut_7 = 14'b11000101011110;
9'd177   : cube_lut_7 = 14'b11000101011111;
9'd178   : cube_lut_7 = 14'b11000101100000;
9'd179   : cube_lut_7 = 14'b11000101100001;
9'd180   : cube_lut_7 = 14'b11000101100010;
9'd181   : cube_lut_7 = 14'b11000101100011;
9'd182   : cube_lut_7 = 14'b11000101100100;
9'd183   : cube_lut_7 = 14'b11000101100110;
9'd184   : cube_lut_7 = 14'b11000101100111;
9'd185   : cube_lut_7 = 14'b11000101101000;
9'd186   : cube_lut_7 = 14'b11000101101001;
9'd187   : cube_lut_7 = 14'b11000101101010;
9'd188   : cube_lut_7 = 14'b11000101101011;
9'd189   : cube_lut_7 = 14'b11000101101100;
9'd190   : cube_lut_7 = 14'b11000101101101;
9'd191   : cube_lut_7 = 14'b11000101101111;
9'd192   : cube_lut_7 = 14'b11000101110000;
9'd193   : cube_lut_7 = 14'b11000101110001;
9'd194   : cube_lut_7 = 14'b11000101110010;
9'd195   : cube_lut_7 = 14'b11000101110011;
9'd196   : cube_lut_7 = 14'b11000101110100;
9'd197   : cube_lut_7 = 14'b11000101110101;
9'd198   : cube_lut_7 = 14'b11000101110110;
9'd199   : cube_lut_7 = 14'b11000101110111;
9'd200   : cube_lut_7 = 14'b11000101111001;
9'd201   : cube_lut_7 = 14'b11000101111010;
9'd202   : cube_lut_7 = 14'b11000101111011;
9'd203   : cube_lut_7 = 14'b11000101111100;
9'd204   : cube_lut_7 = 14'b11000101111101;
9'd205   : cube_lut_7 = 14'b11000101111110;
9'd206   : cube_lut_7 = 14'b11000101111111;
9'd207   : cube_lut_7 = 14'b11000110000000;
9'd208   : cube_lut_7 = 14'b11000110000001;
9'd209   : cube_lut_7 = 14'b11000110000011;
9'd210   : cube_lut_7 = 14'b11000110000100;
9'd211   : cube_lut_7 = 14'b11000110000101;
9'd212   : cube_lut_7 = 14'b11000110000110;
9'd213   : cube_lut_7 = 14'b11000110000111;
9'd214   : cube_lut_7 = 14'b11000110001000;
9'd215   : cube_lut_7 = 14'b11000110001001;
9'd216   : cube_lut_7 = 14'b11000110001010;
9'd217   : cube_lut_7 = 14'b11000110001011;
9'd218   : cube_lut_7 = 14'b11000110001101;
9'd219   : cube_lut_7 = 14'b11000110001110;
9'd220   : cube_lut_7 = 14'b11000110001111;
9'd221   : cube_lut_7 = 14'b11000110010000;
9'd222   : cube_lut_7 = 14'b11000110010001;
9'd223   : cube_lut_7 = 14'b11000110010010;
9'd224   : cube_lut_7 = 14'b11000110010011;
9'd225   : cube_lut_7 = 14'b11000110010100;
9'd226   : cube_lut_7 = 14'b11000110010101;
9'd227   : cube_lut_7 = 14'b11000110010111;
9'd228   : cube_lut_7 = 14'b11000110011000;
9'd229   : cube_lut_7 = 14'b11000110011001;
9'd230   : cube_lut_7 = 14'b11000110011010;
9'd231   : cube_lut_7 = 14'b11000110011011;
9'd232   : cube_lut_7 = 14'b11000110011100;
9'd233   : cube_lut_7 = 14'b11000110011101;
9'd234   : cube_lut_7 = 14'b11000110011110;
9'd235   : cube_lut_7 = 14'b11000110011111;
9'd236   : cube_lut_7 = 14'b11000110100001;
9'd237   : cube_lut_7 = 14'b11000110100010;
9'd238   : cube_lut_7 = 14'b11000110100011;
9'd239   : cube_lut_7 = 14'b11000110100100;
9'd240   : cube_lut_7 = 14'b11000110100101;
9'd241   : cube_lut_7 = 14'b11000110100110;
9'd242   : cube_lut_7 = 14'b11000110100111;
9'd243   : cube_lut_7 = 14'b11000110101000;
9'd244   : cube_lut_7 = 14'b11000110101001;
9'd245   : cube_lut_7 = 14'b11000110101011;
9'd246   : cube_lut_7 = 14'b11000110101100;
9'd247   : cube_lut_7 = 14'b11000110101101;
9'd248   : cube_lut_7 = 14'b11000110101110;
9'd249   : cube_lut_7 = 14'b11000110101111;
9'd250   : cube_lut_7 = 14'b11000110110000;
9'd251   : cube_lut_7 = 14'b11000110110001;
9'd252   : cube_lut_7 = 14'b11000110110010;
9'd253   : cube_lut_7 = 14'b11000110110011;
9'd254   : cube_lut_7 = 14'b11000110110101;
9'd255   : cube_lut_7 = 14'b11000110110110;
9'd256   : cube_lut_7 = 14'b11000110110111;
9'd257   : cube_lut_7 = 14'b11000110111000;
9'd258   : cube_lut_7 = 14'b11000110111001;
9'd259   : cube_lut_7 = 14'b11000110111010;
9'd260   : cube_lut_7 = 14'b11000110111011;
9'd261   : cube_lut_7 = 14'b11000110111100;
9'd262   : cube_lut_7 = 14'b11000110111101;
9'd263   : cube_lut_7 = 14'b11000110111110;
9'd264   : cube_lut_7 = 14'b11000111000000;
9'd265   : cube_lut_7 = 14'b11000111000001;
9'd266   : cube_lut_7 = 14'b11000111000010;
9'd267   : cube_lut_7 = 14'b11000111000011;
9'd268   : cube_lut_7 = 14'b11000111000100;
9'd269   : cube_lut_7 = 14'b11000111000101;
9'd270   : cube_lut_7 = 14'b11000111000110;
9'd271   : cube_lut_7 = 14'b11000111000111;
9'd272   : cube_lut_7 = 14'b11000111001000;
9'd273   : cube_lut_7 = 14'b11000111001001;
9'd274   : cube_lut_7 = 14'b11000111001011;
9'd275   : cube_lut_7 = 14'b11000111001100;
9'd276   : cube_lut_7 = 14'b11000111001101;
9'd277   : cube_lut_7 = 14'b11000111001110;
9'd278   : cube_lut_7 = 14'b11000111001111;
9'd279   : cube_lut_7 = 14'b11000111010000;
9'd280   : cube_lut_7 = 14'b11000111010001;
9'd281   : cube_lut_7 = 14'b11000111010010;
9'd282   : cube_lut_7 = 14'b11000111010011;
9'd283   : cube_lut_7 = 14'b11000111010100;
9'd284   : cube_lut_7 = 14'b11000111010110;
9'd285   : cube_lut_7 = 14'b11000111010111;
9'd286   : cube_lut_7 = 14'b11000111011000;
9'd287   : cube_lut_7 = 14'b11000111011001;
9'd288   : cube_lut_7 = 14'b11000111011010;
9'd289   : cube_lut_7 = 14'b11000111011011;
9'd290   : cube_lut_7 = 14'b11000111011100;
9'd291   : cube_lut_7 = 14'b11000111011101;
9'd292   : cube_lut_7 = 14'b11000111011110;
9'd293   : cube_lut_7 = 14'b11000111011111;
9'd294   : cube_lut_7 = 14'b11000111100001;
9'd295   : cube_lut_7 = 14'b11000111100010;
9'd296   : cube_lut_7 = 14'b11000111100011;
9'd297   : cube_lut_7 = 14'b11000111100100;
9'd298   : cube_lut_7 = 14'b11000111100101;
9'd299   : cube_lut_7 = 14'b11000111100110;
9'd300   : cube_lut_7 = 14'b11000111100111;
9'd301   : cube_lut_7 = 14'b11000111101000;
9'd302   : cube_lut_7 = 14'b11000111101001;
9'd303   : cube_lut_7 = 14'b11000111101010;
9'd304   : cube_lut_7 = 14'b11000111101100;
9'd305   : cube_lut_7 = 14'b11000111101101;
9'd306   : cube_lut_7 = 14'b11000111101110;
9'd307   : cube_lut_7 = 14'b11000111101111;
9'd308   : cube_lut_7 = 14'b11000111110000;
9'd309   : cube_lut_7 = 14'b11000111110001;
9'd310   : cube_lut_7 = 14'b11000111110010;
9'd311   : cube_lut_7 = 14'b11000111110011;
9'd312   : cube_lut_7 = 14'b11000111110100;
9'd313   : cube_lut_7 = 14'b11000111110101;
9'd314   : cube_lut_7 = 14'b11000111110110;
9'd315   : cube_lut_7 = 14'b11000111111000;
9'd316   : cube_lut_7 = 14'b11000111111001;
9'd317   : cube_lut_7 = 14'b11000111111010;
9'd318   : cube_lut_7 = 14'b11000111111011;
9'd319   : cube_lut_7 = 14'b11000111111100;
9'd320   : cube_lut_7 = 14'b11000111111101;
9'd321   : cube_lut_7 = 14'b11000111111110;
9'd322   : cube_lut_7 = 14'b11000111111111;
9'd323   : cube_lut_7 = 14'b11001000000000;
9'd324   : cube_lut_7 = 14'b11001000000001;
9'd325   : cube_lut_7 = 14'b11001000000011;
9'd326   : cube_lut_7 = 14'b11001000000100;
9'd327   : cube_lut_7 = 14'b11001000000101;
9'd328   : cube_lut_7 = 14'b11001000000110;
9'd329   : cube_lut_7 = 14'b11001000000111;
9'd330   : cube_lut_7 = 14'b11001000001000;
9'd331   : cube_lut_7 = 14'b11001000001001;
9'd332   : cube_lut_7 = 14'b11001000001010;
9'd333   : cube_lut_7 = 14'b11001000001011;
9'd334   : cube_lut_7 = 14'b11001000001100;
9'd335   : cube_lut_7 = 14'b11001000001101;
9'd336   : cube_lut_7 = 14'b11001000001111;
9'd337   : cube_lut_7 = 14'b11001000010000;
9'd338   : cube_lut_7 = 14'b11001000010001;
9'd339   : cube_lut_7 = 14'b11001000010010;
9'd340   : cube_lut_7 = 14'b11001000010011;
9'd341   : cube_lut_7 = 14'b11001000010100;
9'd342   : cube_lut_7 = 14'b11001000010101;
9'd343   : cube_lut_7 = 14'b11001000010110;
9'd344   : cube_lut_7 = 14'b11001000010111;
9'd345   : cube_lut_7 = 14'b11001000011000;
9'd346   : cube_lut_7 = 14'b11001000011001;
9'd347   : cube_lut_7 = 14'b11001000011010;
9'd348   : cube_lut_7 = 14'b11001000011100;
9'd349   : cube_lut_7 = 14'b11001000011101;
9'd350   : cube_lut_7 = 14'b11001000011110;
9'd351   : cube_lut_7 = 14'b11001000011111;
9'd352   : cube_lut_7 = 14'b11001000100000;
9'd353   : cube_lut_7 = 14'b11001000100001;
9'd354   : cube_lut_7 = 14'b11001000100010;
9'd355   : cube_lut_7 = 14'b11001000100011;
9'd356   : cube_lut_7 = 14'b11001000100100;
9'd357   : cube_lut_7 = 14'b11001000100101;
9'd358   : cube_lut_7 = 14'b11001000100110;
9'd359   : cube_lut_7 = 14'b11001000101000;
9'd360   : cube_lut_7 = 14'b11001000101001;
9'd361   : cube_lut_7 = 14'b11001000101010;
9'd362   : cube_lut_7 = 14'b11001000101011;
9'd363   : cube_lut_7 = 14'b11001000101100;
9'd364   : cube_lut_7 = 14'b11001000101101;
9'd365   : cube_lut_7 = 14'b11001000101110;
9'd366   : cube_lut_7 = 14'b11001000101111;
9'd367   : cube_lut_7 = 14'b11001000110000;
9'd368   : cube_lut_7 = 14'b11001000110001;
9'd369   : cube_lut_7 = 14'b11001000110010;
9'd370   : cube_lut_7 = 14'b11001000110011;
9'd371   : cube_lut_7 = 14'b11001000110101;
9'd372   : cube_lut_7 = 14'b11001000110110;
9'd373   : cube_lut_7 = 14'b11001000110111;
9'd374   : cube_lut_7 = 14'b11001000111000;
9'd375   : cube_lut_7 = 14'b11001000111001;
9'd376   : cube_lut_7 = 14'b11001000111010;
9'd377   : cube_lut_7 = 14'b11001000111011;
9'd378   : cube_lut_7 = 14'b11001000111100;
9'd379   : cube_lut_7 = 14'b11001000111101;
9'd380   : cube_lut_7 = 14'b11001000111110;
9'd381   : cube_lut_7 = 14'b11001000111111;
9'd382   : cube_lut_7 = 14'b11001001000000;
9'd383   : cube_lut_7 = 14'b11001001000010;
9'd384   : cube_lut_7 = 14'b11001001000011;
9'd385   : cube_lut_7 = 14'b11001001000100;
9'd386   : cube_lut_7 = 14'b11001001000101;
9'd387   : cube_lut_7 = 14'b11001001000110;
9'd388   : cube_lut_7 = 14'b11001001000111;
9'd389   : cube_lut_7 = 14'b11001001001000;
9'd390   : cube_lut_7 = 14'b11001001001001;
9'd391   : cube_lut_7 = 14'b11001001001010;
9'd392   : cube_lut_7 = 14'b11001001001011;
9'd393   : cube_lut_7 = 14'b11001001001100;
9'd394   : cube_lut_7 = 14'b11001001001101;
9'd395   : cube_lut_7 = 14'b11001001001110;
9'd396   : cube_lut_7 = 14'b11001001010000;
9'd397   : cube_lut_7 = 14'b11001001010001;
9'd398   : cube_lut_7 = 14'b11001001010010;
9'd399   : cube_lut_7 = 14'b11001001010011;
9'd400   : cube_lut_7 = 14'b11001001010100;
9'd401   : cube_lut_7 = 14'b11001001010101;
9'd402   : cube_lut_7 = 14'b11001001010110;
9'd403   : cube_lut_7 = 14'b11001001010111;
9'd404   : cube_lut_7 = 14'b11001001011000;
9'd405   : cube_lut_7 = 14'b11001001011001;
9'd406   : cube_lut_7 = 14'b11001001011010;
9'd407   : cube_lut_7 = 14'b11001001011011;
9'd408   : cube_lut_7 = 14'b11001001011100;
9'd409   : cube_lut_7 = 14'b11001001011110;
9'd410   : cube_lut_7 = 14'b11001001011111;
9'd411   : cube_lut_7 = 14'b11001001100000;
9'd412   : cube_lut_7 = 14'b11001001100001;
9'd413   : cube_lut_7 = 14'b11001001100010;
9'd414   : cube_lut_7 = 14'b11001001100011;
9'd415   : cube_lut_7 = 14'b11001001100100;
9'd416   : cube_lut_7 = 14'b11001001100101;
9'd417   : cube_lut_7 = 14'b11001001100110;
9'd418   : cube_lut_7 = 14'b11001001100111;
9'd419   : cube_lut_7 = 14'b11001001101000;
9'd420   : cube_lut_7 = 14'b11001001101001;
9'd421   : cube_lut_7 = 14'b11001001101010;
9'd422   : cube_lut_7 = 14'b11001001101100;
9'd423   : cube_lut_7 = 14'b11001001101101;
9'd424   : cube_lut_7 = 14'b11001001101110;
9'd425   : cube_lut_7 = 14'b11001001101111;
9'd426   : cube_lut_7 = 14'b11001001110000;
9'd427   : cube_lut_7 = 14'b11001001110001;
9'd428   : cube_lut_7 = 14'b11001001110010;
9'd429   : cube_lut_7 = 14'b11001001110011;
9'd430   : cube_lut_7 = 14'b11001001110100;
9'd431   : cube_lut_7 = 14'b11001001110101;
9'd432   : cube_lut_7 = 14'b11001001110110;
9'd433   : cube_lut_7 = 14'b11001001110111;
9'd434   : cube_lut_7 = 14'b11001001111000;
9'd435   : cube_lut_7 = 14'b11001001111001;
9'd436   : cube_lut_7 = 14'b11001001111011;
9'd437   : cube_lut_7 = 14'b11001001111100;
9'd438   : cube_lut_7 = 14'b11001001111101;
9'd439   : cube_lut_7 = 14'b11001001111110;
9'd440   : cube_lut_7 = 14'b11001001111111;
9'd441   : cube_lut_7 = 14'b11001010000000;
9'd442   : cube_lut_7 = 14'b11001010000001;
9'd443   : cube_lut_7 = 14'b11001010000010;
9'd444   : cube_lut_7 = 14'b11001010000011;
9'd445   : cube_lut_7 = 14'b11001010000100;
9'd446   : cube_lut_7 = 14'b11001010000101;
9'd447   : cube_lut_7 = 14'b11001010000110;
9'd448   : cube_lut_7 = 14'b11001010000111;
9'd449   : cube_lut_7 = 14'b11001010001000;
9'd450   : cube_lut_7 = 14'b11001010001010;
9'd451   : cube_lut_7 = 14'b11001010001011;
9'd452   : cube_lut_7 = 14'b11001010001100;
9'd453   : cube_lut_7 = 14'b11001010001101;
9'd454   : cube_lut_7 = 14'b11001010001110;
9'd455   : cube_lut_7 = 14'b11001010001111;
9'd456   : cube_lut_7 = 14'b11001010010000;
9'd457   : cube_lut_7 = 14'b11001010010001;
9'd458   : cube_lut_7 = 14'b11001010010010;
9'd459   : cube_lut_7 = 14'b11001010010011;
9'd460   : cube_lut_7 = 14'b11001010010100;
9'd461   : cube_lut_7 = 14'b11001010010101;
9'd462   : cube_lut_7 = 14'b11001010010110;
9'd463   : cube_lut_7 = 14'b11001010010111;
9'd464   : cube_lut_7 = 14'b11001010011000;
9'd465   : cube_lut_7 = 14'b11001010011010;
9'd466   : cube_lut_7 = 14'b11001010011011;
9'd467   : cube_lut_7 = 14'b11001010011100;
9'd468   : cube_lut_7 = 14'b11001010011101;
9'd469   : cube_lut_7 = 14'b11001010011110;
9'd470   : cube_lut_7 = 14'b11001010011111;
9'd471   : cube_lut_7 = 14'b11001010100000;
9'd472   : cube_lut_7 = 14'b11001010100001;
9'd473   : cube_lut_7 = 14'b11001010100010;
9'd474   : cube_lut_7 = 14'b11001010100011;
9'd475   : cube_lut_7 = 14'b11001010100100;
9'd476   : cube_lut_7 = 14'b11001010100101;
9'd477   : cube_lut_7 = 14'b11001010100110;
9'd478   : cube_lut_7 = 14'b11001010100111;
9'd479   : cube_lut_7 = 14'b11001010101000;
9'd480   : cube_lut_7 = 14'b11001010101010;
9'd481   : cube_lut_7 = 14'b11001010101011;
9'd482   : cube_lut_7 = 14'b11001010101100;
9'd483   : cube_lut_7 = 14'b11001010101101;
9'd484   : cube_lut_7 = 14'b11001010101110;
9'd485   : cube_lut_7 = 14'b11001010101111;
9'd486   : cube_lut_7 = 14'b11001010110000;
9'd487   : cube_lut_7 = 14'b11001010110001;
9'd488   : cube_lut_7 = 14'b11001010110010;
9'd489   : cube_lut_7 = 14'b11001010110011;
9'd490   : cube_lut_7 = 14'b11001010110100;
9'd491   : cube_lut_7 = 14'b11001010110101;
9'd492   : cube_lut_7 = 14'b11001010110110;
9'd493   : cube_lut_7 = 14'b11001010110111;
9'd494   : cube_lut_7 = 14'b11001010111000;
9'd495   : cube_lut_7 = 14'b11001010111001;
9'd496   : cube_lut_7 = 14'b11001010111011;
9'd497   : cube_lut_7 = 14'b11001010111100;
9'd498   : cube_lut_7 = 14'b11001010111101;
9'd499   : cube_lut_7 = 14'b11001010111110;
9'd500   : cube_lut_7 = 14'b11001010111111;
9'd501   : cube_lut_7 = 14'b11001011000000;
9'd502   : cube_lut_7 = 14'b11001011000001;
9'd503   : cube_lut_7 = 14'b11001011000010;
9'd504   : cube_lut_7 = 14'b11001011000011;
9'd505   : cube_lut_7 = 14'b11001011000100;
9'd506   : cube_lut_7 = 14'b11001011000101;
9'd507   : cube_lut_7 = 14'b11001011000110;
9'd508   : cube_lut_7 = 14'b11001011000111;
9'd509   : cube_lut_7 = 14'b11001011001000;
9'd510   : cube_lut_7 = 14'b11001011001001;
9'd511   : cube_lut_7 = 14'b11001011001010;

    endcase
end

//----------------------------------------------//
// Module Instance                              //
//----------------------------------------------//

always@(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        o_data      <= 0;
        o_prcis_idx <= 0;
    end
    else begin
        o_data      <= o_data_nxt;
        o_prcis_idx <= o_prcis_idx_nxt;
    end
end

endmodule

