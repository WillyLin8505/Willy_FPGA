parameter SSR_PX_FMT   = "RGB16";
parameter MON_PX_FMT   = "RGB8";
parameter GENERATE_SEL = 1;
parameter OUT_TYPE     = "YCBCR";
parameter           YCBCR_POS               = 0;
parameter           CIIW_RY                 = 8; //rgb   integer precision
parameter           CIPW_RY                 = 0; //rgb   point   precision 
parameter           COIW_RY                 = 8; //ycbcr integer precision 
parameter           COPW_RY                 = 4; //ycbcr point   precision 
parameter           CIIW_YL                 = 8; //ycbcr integer precision 
parameter           CIPW_YL                 = 4; //ycbcr point   precision 
parameter           COIW_YL                 = 8; //lms   integer precision 
parameter           COPW_YL                 = 4; //lms   point   precision 
parameter           CIIW_LK                 = 8; //lms   integer precision 
parameter           CIPW_LK                 = 4; //lms   point   precision
parameter           COIW_L_LK               = 0; //l     inetger precision 
parameter           COPW_L_LK               = 15;//l     point   precision
parameter           COIW_AB_LK              = 1; //ab    inetger precision 
parameter           COPW_AB_LK              = 13;//ab    point   precision
parameter           CIIW_KL                 = 0; //l     inetger precision 
parameter           CIPW_KL                 = 15;//l     point   precision
parameter           CIIW_KAB                = 1; //ab    inetger precision 
parameter           CIPW_KAB                = 13;//ab    point   precision
parameter           CIW_LMS                 = 0; //lms   integer precision 
parameter           CPW_LMS                 = 15;//lms   point   precision
parameter           CIW_STG_1_KL            = 0; //mul stage 1   precision 
parameter           CPW_STG_1_KL            = 14;//mul stage 2   precision 
parameter           COIW_KL                 = 8; //cube  integer precision 
parameter           COPW_KL                 = 6; //cube  point   precision
parameter           CIIW_LR                 = 8; //cube  integer precision 
parameter           CIPW_LR                 = 6; //cube  point   precision
parameter           COIW_LR                 = 8; //rgb   integer precision 
parameter           COPW_LR                 = 0; //rgb   point   precision 
parameter           COIW_LY                 = 8; //ycbcr integer precision 
parameter           COPW_LY                 = 4; //ycbcr point   precision 
