parameter  SSR_PX_FMT       = "RGB10";
parameter  DBUF_DW          = 10;
parameter  RAW_CIIW         = DBUF_DW;
parameter  RAW_CIPW         = 0;
parameter  DPC_NUM          = 2;
parameter  INS_CIW          = DBUF_DW*2;
parameter  ALG_LVL          = "LVL_0";
parameter  ALG_MODE         = "SDPC";
parameter  IMG_HSZ          = 1928;
parameter  IMG_VSZ          = 1080;
parameter ODATA_FREQ       = 0;
parameter BUF_PIXEL_DLY    = 0;
parameter BUF_LINE_DLY     = 0;
parameter MEM_TYPE         = "1PSRAM";
parameter SRAM_SEL         = 2;
parameter MEM_NAME         = (SRAM_SEL == 1) ? "asic_sram_sp240x160" : "M31HDSP100PL040P_488X1X80CM4";
parameter SRAM_NUM         = (SRAM_SEL == 1) ? 1 : 2;
