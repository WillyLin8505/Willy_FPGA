    parameter DBUF_DW      = 8;
    parameter DBUF_DEP     = 1920;
    parameter KRNV_SZ      = 5;                     // vertical kernel size
    parameter KRNH_SZ      = 5;                     // horizontial kernel size
    parameter ODATA_RNG    = 3;                     // output data range //cannot set to 1 
    parameter ODATA_FREQ   = 0;                     // output data frequence : 0:every 1 cycle change output data 
    parameter TOP_PAD      = 2;                     // top padding line number 
    parameter BTM_PAD      = 2;                     // bottom padding line number 
    parameter FR_PAD       = 1;                     // front padding number 
    parameter BK_PAD       = 1;                     // back padding number 
    parameter PAD_MODE     = 0;                     // 0:for duplicate padding 
    parameter BUF_PIXEL_DLY    = 0;
    parameter BUF_LINE_DLY     = 0;
    parameter SEN_PIXEL_DLY    = 1;
