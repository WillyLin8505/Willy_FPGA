parameter SSR_PX_FMT  = "RGB16";
parameter MON_PX_FMT= "RGB14";
parameter  IMG_HSZ= 32768;
parameter  IMG_VSZ= 1;
parameter  CIIW= 0;
parameter  CIPW= 15;
parameter  COIW= 0;
parameter  COPW= 13;
parameter  SEL_CURVE = "OK_L";
parameter  CIW= CIIW + CIPW;
parameter  COW=  COIW + COPW;
parameter  LUT_MAP_WTH =  (SEL_CURVE== "REFI_L") ? 11 : (SEL_CURVE== "REFI_C") ? 8  : 13;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_0= 0;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_1= 697;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_2= 973;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_3= 1232;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_4= 1718;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_5= 2176;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_6= 2598;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_7= 2972;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_8= 3311;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_9= 3625;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_10= 3918;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_11= 4194;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_12= 4457;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_13= 4708;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_14= 4948;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_15= 5180;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_16= 5620;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_17= 6034;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_18= 6426;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_19= 6800;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_20= 7158;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_21= 7502;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_22= 7804;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_23= 8045;
parameter  [LUT_MAP_WTH-1:0] Y_DATA_24= 8191;
