parameter SSR_PX_FMT    ="RGB8";
parameter YCBCR_COIW    =8;
parameter YCBCR_COPW    =4;
parameter LINE_BUF_COIW =YCBCR_COIW;
parameter LINE_BUF_COPW =YCBCR_COPW;
parameter BIL_FTR_COIW  =LINE_BUF_COIW;
parameter BIL_FTR_COPW  =LINE_BUF_COPW;
parameter DUF_DEP       =1920;
parameter IMG_HSZ       =1920;
parameter IMG_VSZ       =1080; 
parameter YCBCR_POS     =0;
parameter KRNV_SZ       =5;                   // vertical kernel size
parameter KRNH_SZ       =5;                    // horizontial kernel size 
parameter ODATA_RNG     =5;                   // output data range //cannot set to 1 
parameter ODATA_FREQ    =0;                    // output data frequence : 0:every 1 cycle change output data 
parameter TOP_PAD       =2;                    // top padding line number 
parameter BTM_PAD       =2;                  // bottom padding line number 
parameter FR_PAD        =2;                     // front padding number  
parameter BK_PAD        =2;                      // back padding number 
parameter PAD_MODE      =0;                  // 0:for duplicate padding  1:raw data padding 
parameter SIGN_EN      = 1;
