// +FHDR -----------------------------------------------------------------------
// Copyright (c) Silicon Optronics. Inc. 2022
//
// File Name:           ip_cube_lut_12_14_ver2.v
// Author:              1.Willy Lin
//                      2.Martin Chen
//                      3.Humphrey Lin
// Version:             1.0
// Last Modified On:    2023/1/3
//
// File Description:    cube root lut
// Abbreviations:
// File precision  :    input  : 0.12
//                      output : 0.14

// Consuming time :     1T
// -FHDR -----------------------------------------------------------------------

module ip_cube_lut_12_14_ver2
(
//----------------------------------------------//
// Output declaration                           //
//----------------------------------------------//
    output reg [13:0] o_data,

//----------------------------------------------//
// Input declaration                            //
//----------------------------------------------//
    input      [11:0] i_data,
    input             clk,
    input             rst_n
);

//----------------------------------------------//
// Local Parameter                              //
//----------------------------------------------//

//----------------------------------------------//
// Register & Wire declaration                  //
//----------------------------------------------//
wire        decode_0;
wire        decode_1;
wire        decode_2;
wire        decode_3;

wire [13:0] com_lut;

reg  [13:0] cube_lut_0;
reg  [13:0] cube_lut_1;
reg  [13:0] cube_lut_2;
reg  [13:0] cube_lut_3;

//output port
wire [13:0] o_data_nxt;

//----------------------------------------------//
// Code Descriptions                            //
//----------------------------------------------//
//find region
assign decode_0 = i_data[11:10] == 2'b00;
assign decode_1 = i_data[11:10] == 2'b01;
assign decode_2 = i_data[11:10] == 2'b10;
assign decode_3 = i_data[11:10] == 2'b11;

assign com_lut = ({14{decode_0}} & cube_lut_0) |
                 ({14{decode_1}} & cube_lut_1) |
                 ({14{decode_2}} & cube_lut_2) |
                 ({14{decode_3}} & cube_lut_3);

assign o_data_nxt = com_lut;

always@* begin
    
    cube_lut_0 = 0;
    
    case(i_data[9:0])
        10'd0   : cube_lut_0    = 14'b00000000000000;
        10'd1   : cube_lut_0    = 14'b00010000000000;
        10'd2   : cube_lut_0    = 14'b00010100001010;
        10'd3   : cube_lut_0    = 14'b00010111000100;
        10'd4   : cube_lut_0    = 14'b00011001011001;
        10'd5   : cube_lut_0    = 14'b00011011010111;
        10'd6   : cube_lut_0    = 14'b00011101000100;
        10'd7   : cube_lut_0    = 14'b00011110100110;
        10'd8   : cube_lut_0    = 14'b00100000000000;
        10'd9   : cube_lut_0    = 14'b00100001010010;
        10'd10   : cube_lut_0   = 14'b00100010011110;
        10'd11   : cube_lut_0   = 14'b00100011100101;
        10'd12   : cube_lut_0   = 14'b00100100101000;
        10'd13   : cube_lut_0   = 14'b00100101100111;
        10'd14   : cube_lut_0   = 14'b00100110100011;
        10'd15   : cube_lut_0   = 14'b00100111011101;
        10'd16   : cube_lut_0   = 14'b00101000010100;
        10'd17   : cube_lut_0   = 14'b00101001001000;
        10'd18   : cube_lut_0   = 14'b00101001111011;
        10'd19   : cube_lut_0   = 14'b00101010101100;
        10'd20   : cube_lut_0   = 14'b00101011011011;
        10'd21   : cube_lut_0   = 14'b00101100001001;
        10'd22   : cube_lut_0   = 14'b00101100110101;
        10'd23   : cube_lut_0   = 14'b00101101100000;
        10'd24   : cube_lut_0   = 14'b00101110001001;
        10'd25   : cube_lut_0   = 14'b00101110110010;
        10'd26   : cube_lut_0   = 14'b00101111011001;
        10'd27   : cube_lut_0   = 14'b00110000000000;
        10'd28   : cube_lut_0   = 14'b00110000100101;
        10'd29   : cube_lut_0   = 14'b00110001001010;
        10'd30   : cube_lut_0   = 14'b00110001101101;
        10'd31   : cube_lut_0   = 14'b00110010010000;
        10'd32   : cube_lut_0   = 14'b00110010110010;
        10'd33   : cube_lut_0   = 14'b00110011010100;
        10'd34   : cube_lut_0   = 14'b00110011110101;
        10'd35   : cube_lut_0   = 14'b00110100010101;
        10'd36   : cube_lut_0   = 14'b00110100110101;
        10'd37   : cube_lut_0   = 14'b00110101010100;
        10'd38   : cube_lut_0   = 14'b00110101110010;
        10'd39   : cube_lut_0   = 14'b00110110010000;
        10'd40   : cube_lut_0   = 14'b00110110101110;
        10'd41   : cube_lut_0   = 14'b00110111001010;
        10'd42   : cube_lut_0   = 14'b00110111100111;
        10'd43   : cube_lut_0   = 14'b00111000000011;
        10'd44   : cube_lut_0   = 14'b00111000011111;
        10'd45   : cube_lut_0   = 14'b00111000111010;
        10'd46   : cube_lut_0   = 14'b00111001010101;
        10'd47   : cube_lut_0   = 14'b00111001101111;
        10'd48   : cube_lut_0   = 14'b00111010001001;
        10'd49   : cube_lut_0   = 14'b00111010100011;
        10'd50   : cube_lut_0   = 14'b00111010111100;
        10'd51   : cube_lut_0   = 14'b00111011010101;
        10'd52   : cube_lut_0   = 14'b00111011101110;
        10'd53   : cube_lut_0   = 14'b00111100000110;
        10'd54   : cube_lut_0   = 14'b00111100011110;
        10'd55   : cube_lut_0   = 14'b00111100110110;
        10'd56   : cube_lut_0   = 14'b00111101001101;
        10'd57   : cube_lut_0   = 14'b00111101100100;
        10'd58   : cube_lut_0   = 14'b00111101111011;
        10'd59   : cube_lut_0   = 14'b00111110010010;
        10'd60   : cube_lut_0   = 14'b00111110101000;
        10'd61   : cube_lut_0   = 14'b00111110111110;
        10'd62   : cube_lut_0   = 14'b00111111010100;
        10'd63   : cube_lut_0   = 14'b00111111101010;
        10'd64   : cube_lut_0   = 14'b01000000000000;
        10'd65   : cube_lut_0   = 14'b01000000010101;
        10'd66   : cube_lut_0   = 14'b01000000101010;
        10'd67   : cube_lut_0   = 14'b01000000111111;
        10'd68   : cube_lut_0   = 14'b01000001010011;
        10'd69   : cube_lut_0   = 14'b01000001101000;
        10'd70   : cube_lut_0   = 14'b01000001111100;
        10'd71   : cube_lut_0   = 14'b01000010010000;
        10'd72   : cube_lut_0   = 14'b01000010100100;
        10'd73   : cube_lut_0   = 14'b01000010110111;
        10'd74   : cube_lut_0   = 14'b01000011001011;
        10'd75   : cube_lut_0   = 14'b01000011011110;
        10'd76   : cube_lut_0   = 14'b01000011110001;
        10'd77   : cube_lut_0   = 14'b01000100000100;
        10'd78   : cube_lut_0   = 14'b01000100010111;
        10'd79   : cube_lut_0   = 14'b01000100101001;
        10'd80   : cube_lut_0   = 14'b01000100111100;
        10'd81   : cube_lut_0   = 14'b01000101001110;
        10'd82   : cube_lut_0   = 14'b01000101100000;
        10'd83   : cube_lut_0   = 14'b01000101110010;
        10'd84   : cube_lut_0   = 14'b01000110000100;
        10'd85   : cube_lut_0   = 14'b01000110010110;
        10'd86   : cube_lut_0   = 14'b01000110100111;
        10'd87   : cube_lut_0   = 14'b01000110111001;
        10'd88   : cube_lut_0   = 14'b01000111001010;
        10'd89   : cube_lut_0   = 14'b01000111011011;
        10'd90   : cube_lut_0   = 14'b01000111101100;
        10'd91   : cube_lut_0   = 14'b01000111111101;
        10'd92   : cube_lut_0   = 14'b01001000001110;
        10'd93   : cube_lut_0   = 14'b01001000011111;
        10'd94   : cube_lut_0   = 14'b01001000101111;
        10'd95   : cube_lut_0   = 14'b01001001000000;
        10'd96   : cube_lut_0   = 14'b01001001010000;
        10'd97   : cube_lut_0   = 14'b01001001100000;
        10'd98   : cube_lut_0   = 14'b01001001110001;
        10'd99   : cube_lut_0   = 14'b01001010000001;
        10'd100   : cube_lut_0  = 14'b01001010010000;
        10'd101   : cube_lut_0  = 14'b01001010100000;
        10'd102   : cube_lut_0  = 14'b01001010110000;
        10'd103   : cube_lut_0  = 14'b01001011000000;
        10'd104   : cube_lut_0  = 14'b01001011001111;
        10'd105   : cube_lut_0  = 14'b01001011011110;
        10'd106   : cube_lut_0  = 14'b01001011101110;
        10'd107   : cube_lut_0  = 14'b01001011111101;
        10'd108   : cube_lut_0  = 14'b01001100001100;
        10'd109   : cube_lut_0  = 14'b01001100011011;
        10'd110   : cube_lut_0  = 14'b01001100101010;
        10'd111   : cube_lut_0  = 14'b01001100111001;
        10'd112   : cube_lut_0  = 14'b01001101000111;
        10'd113   : cube_lut_0  = 14'b01001101010110;
        10'd114   : cube_lut_0  = 14'b01001101100101;
        10'd115   : cube_lut_0  = 14'b01001101110011;
        10'd116   : cube_lut_0  = 14'b01001110000010;
        10'd117   : cube_lut_0  = 14'b01001110010000;
        10'd118   : cube_lut_0  = 14'b01001110011110;
        10'd119   : cube_lut_0  = 14'b01001110101100;
        10'd120   : cube_lut_0  = 14'b01001110111010;
        10'd121   : cube_lut_0  = 14'b01001111001000;
        10'd122   : cube_lut_0  = 14'b01001111010110;
        10'd123   : cube_lut_0  = 14'b01001111100100;
        10'd124   : cube_lut_0  = 14'b01001111110010;
        10'd125   : cube_lut_0  = 14'b01010000000000;
        10'd126   : cube_lut_0  = 14'b01010000001101;
        10'd127   : cube_lut_0  = 14'b01010000011011;
        10'd128   : cube_lut_0  = 14'b01010000101000;
        10'd129   : cube_lut_0  = 14'b01010000110110;
        10'd130   : cube_lut_0  = 14'b01010001000011;
        10'd131   : cube_lut_0  = 14'b01010001010000;
        10'd132   : cube_lut_0  = 14'b01010001011101;
        10'd133   : cube_lut_0  = 14'b01010001101010;
        10'd134   : cube_lut_0  = 14'b01010001111000;
        10'd135   : cube_lut_0  = 14'b01010010000101;
        10'd136   : cube_lut_0  = 14'b01010010010001;
        10'd137   : cube_lut_0  = 14'b01010010011110;
        10'd138   : cube_lut_0  = 14'b01010010101011;
        10'd139   : cube_lut_0  = 14'b01010010111000;
        10'd140   : cube_lut_0  = 14'b01010011000101;
        10'd141   : cube_lut_0  = 14'b01010011010001;
        10'd142   : cube_lut_0  = 14'b01010011011110;
        10'd143   : cube_lut_0  = 14'b01010011101010;
        10'd144   : cube_lut_0  = 14'b01010011110111;
        10'd145   : cube_lut_0  = 14'b01010100000011;
        10'd146   : cube_lut_0  = 14'b01010100010000;
        10'd147   : cube_lut_0  = 14'b01010100011100;
        10'd148   : cube_lut_0  = 14'b01010100101000;
        10'd149   : cube_lut_0  = 14'b01010100110100;
        10'd150   : cube_lut_0  = 14'b01010101000000;
        10'd151   : cube_lut_0  = 14'b01010101001100;
        10'd152   : cube_lut_0  = 14'b01010101011000;
        10'd153   : cube_lut_0  = 14'b01010101100100;
        10'd154   : cube_lut_0  = 14'b01010101110000;
        10'd155   : cube_lut_0  = 14'b01010101111100;
        10'd156   : cube_lut_0  = 14'b01010110001000;
        10'd157   : cube_lut_0  = 14'b01010110010100;
        10'd158   : cube_lut_0  = 14'b01010110011111;
        10'd159   : cube_lut_0  = 14'b01010110101011;
        10'd160   : cube_lut_0  = 14'b01010110110111;
        10'd161   : cube_lut_0  = 14'b01010111000010;
        10'd162   : cube_lut_0  = 14'b01010111001110;
        10'd163   : cube_lut_0  = 14'b01010111011001;
        10'd164   : cube_lut_0  = 14'b01010111100101;
        10'd165   : cube_lut_0  = 14'b01010111110000;
        10'd166   : cube_lut_0  = 14'b01010111111011;
        10'd167   : cube_lut_0  = 14'b01011000000111;
        10'd168   : cube_lut_0  = 14'b01011000010010;
        10'd169   : cube_lut_0  = 14'b01011000011101;
        10'd170   : cube_lut_0  = 14'b01011000101000;
        10'd171   : cube_lut_0  = 14'b01011000110011;
        10'd172   : cube_lut_0  = 14'b01011000111110;
        10'd173   : cube_lut_0  = 14'b01011001001001;
        10'd174   : cube_lut_0  = 14'b01011001010100;
        10'd175   : cube_lut_0  = 14'b01011001011111;
        10'd176   : cube_lut_0  = 14'b01011001101010;
        10'd177   : cube_lut_0  = 14'b01011001110101;
        10'd178   : cube_lut_0  = 14'b01011010000000;
        10'd179   : cube_lut_0  = 14'b01011010001010;
        10'd180   : cube_lut_0  = 14'b01011010010101;
        10'd181   : cube_lut_0  = 14'b01011010100000;
        10'd182   : cube_lut_0  = 14'b01011010101011;
        10'd183   : cube_lut_0  = 14'b01011010110101;
        10'd184   : cube_lut_0  = 14'b01011011000000;
        10'd185   : cube_lut_0  = 14'b01011011001010;
        10'd186   : cube_lut_0  = 14'b01011011010101;
        10'd187   : cube_lut_0  = 14'b01011011011111;
        10'd188   : cube_lut_0  = 14'b01011011101010;
        10'd189   : cube_lut_0  = 14'b01011011110100;
        10'd190   : cube_lut_0  = 14'b01011011111110;
        10'd191   : cube_lut_0  = 14'b01011100001001;
        10'd192   : cube_lut_0  = 14'b01011100010011;
        10'd193   : cube_lut_0  = 14'b01011100011101;
        10'd194   : cube_lut_0  = 14'b01011100100111;
        10'd195   : cube_lut_0  = 14'b01011100110010;
        10'd196   : cube_lut_0  = 14'b01011100111100;
        10'd197   : cube_lut_0  = 14'b01011101000110;
        10'd198   : cube_lut_0  = 14'b01011101010000;
        10'd199   : cube_lut_0  = 14'b01011101011010;
        10'd200   : cube_lut_0  = 14'b01011101100100;
        10'd201   : cube_lut_0  = 14'b01011101101110;
        10'd202   : cube_lut_0  = 14'b01011101111000;
        10'd203   : cube_lut_0  = 14'b01011110000010;
        10'd204   : cube_lut_0  = 14'b01011110001100;
        10'd205   : cube_lut_0  = 14'b01011110010101;
        10'd206   : cube_lut_0  = 14'b01011110011111;
        10'd207   : cube_lut_0  = 14'b01011110101001;
        10'd208   : cube_lut_0  = 14'b01011110110011;
        10'd209   : cube_lut_0  = 14'b01011110111100;
        10'd210   : cube_lut_0  = 14'b01011111000110;
        10'd211   : cube_lut_0  = 14'b01011111010000;
        10'd212   : cube_lut_0  = 14'b01011111011001;
        10'd213   : cube_lut_0  = 14'b01011111100011;
        10'd214   : cube_lut_0  = 14'b01011111101100;
        10'd215   : cube_lut_0  = 14'b01011111110110;
        10'd216   : cube_lut_0  = 14'b01100000000000;
        10'd217   : cube_lut_0  = 14'b01100000001001;
        10'd218   : cube_lut_0  = 14'b01100000010010;
        10'd219   : cube_lut_0  = 14'b01100000011100;
        10'd220   : cube_lut_0  = 14'b01100000100101;
        10'd221   : cube_lut_0  = 14'b01100000101111;
        10'd222   : cube_lut_0  = 14'b01100000111000;
        10'd223   : cube_lut_0  = 14'b01100001000001;
        10'd224   : cube_lut_0  = 14'b01100001001010;
        10'd225   : cube_lut_0  = 14'b01100001010100;
        10'd226   : cube_lut_0  = 14'b01100001011101;
        10'd227   : cube_lut_0  = 14'b01100001100110;
        10'd228   : cube_lut_0  = 14'b01100001101111;
        10'd229   : cube_lut_0  = 14'b01100001111000;
        10'd230   : cube_lut_0  = 14'b01100010000001;
        10'd231   : cube_lut_0  = 14'b01100010001011;
        10'd232   : cube_lut_0  = 14'b01100010010100;
        10'd233   : cube_lut_0  = 14'b01100010011101;
        10'd234   : cube_lut_0  = 14'b01100010100110;
        10'd235   : cube_lut_0  = 14'b01100010101111;
        10'd236   : cube_lut_0  = 14'b01100010111000;
        10'd237   : cube_lut_0  = 14'b01100011000000;
        10'd238   : cube_lut_0  = 14'b01100011001001;
        10'd239   : cube_lut_0  = 14'b01100011010010;
        10'd240   : cube_lut_0  = 14'b01100011011011;
        10'd241   : cube_lut_0  = 14'b01100011100100;
        10'd242   : cube_lut_0  = 14'b01100011101101;
        10'd243   : cube_lut_0  = 14'b01100011110110;
        10'd244   : cube_lut_0  = 14'b01100011111110;
        10'd245   : cube_lut_0  = 14'b01100100000111;
        10'd246   : cube_lut_0  = 14'b01100100010000;
        10'd247   : cube_lut_0  = 14'b01100100011000;
        10'd248   : cube_lut_0  = 14'b01100100100001;
        10'd249   : cube_lut_0  = 14'b01100100101010;
        10'd250   : cube_lut_0  = 14'b01100100110010;
        10'd251   : cube_lut_0  = 14'b01100100111011;
        10'd252   : cube_lut_0  = 14'b01100101000011;
        10'd253   : cube_lut_0  = 14'b01100101001100;
        10'd254   : cube_lut_0  = 14'b01100101010101;
        10'd255   : cube_lut_0  = 14'b01100101011101;
        10'd256   : cube_lut_0  = 14'b01100101100101;
        10'd257   : cube_lut_0  = 14'b01100101101110;
        10'd258   : cube_lut_0  = 14'b01100101110110;
        10'd259   : cube_lut_0  = 14'b01100101111111;
        10'd260   : cube_lut_0  = 14'b01100110000111;
        10'd261   : cube_lut_0  = 14'b01100110010000;
        10'd262   : cube_lut_0  = 14'b01100110011000;
        10'd263   : cube_lut_0  = 14'b01100110100000;
        10'd264   : cube_lut_0  = 14'b01100110101001;
        10'd265   : cube_lut_0  = 14'b01100110110001;
        10'd266   : cube_lut_0  = 14'b01100110111001;
        10'd267   : cube_lut_0  = 14'b01100111000001;
        10'd268   : cube_lut_0  = 14'b01100111001010;
        10'd269   : cube_lut_0  = 14'b01100111010010;
        10'd270   : cube_lut_0  = 14'b01100111011010;
        10'd271   : cube_lut_0  = 14'b01100111100010;
        10'd272   : cube_lut_0  = 14'b01100111101010;
        10'd273   : cube_lut_0  = 14'b01100111110010;
        10'd274   : cube_lut_0  = 14'b01100111111010;
        10'd275   : cube_lut_0  = 14'b01101000000011;
        10'd276   : cube_lut_0  = 14'b01101000001011;
        10'd277   : cube_lut_0  = 14'b01101000010011;
        10'd278   : cube_lut_0  = 14'b01101000011011;
        10'd279   : cube_lut_0  = 14'b01101000100011;
        10'd280   : cube_lut_0  = 14'b01101000101011;
        10'd281   : cube_lut_0  = 14'b01101000110011;
        10'd282   : cube_lut_0  = 14'b01101000111011;
        10'd283   : cube_lut_0  = 14'b01101001000010;
        10'd284   : cube_lut_0  = 14'b01101001001010;
        10'd285   : cube_lut_0  = 14'b01101001010010;
        10'd286   : cube_lut_0  = 14'b01101001011010;
        10'd287   : cube_lut_0  = 14'b01101001100010;
        10'd288   : cube_lut_0  = 14'b01101001101010;
        10'd289   : cube_lut_0  = 14'b01101001110010;
        10'd290   : cube_lut_0  = 14'b01101001111001;
        10'd291   : cube_lut_0  = 14'b01101010000001;
        10'd292   : cube_lut_0  = 14'b01101010001001;
        10'd293   : cube_lut_0  = 14'b01101010010001;
        10'd294   : cube_lut_0  = 14'b01101010011000;
        10'd295   : cube_lut_0  = 14'b01101010100000;
        10'd296   : cube_lut_0  = 14'b01101010101000;
        10'd297   : cube_lut_0  = 14'b01101010110000;
        10'd298   : cube_lut_0  = 14'b01101010110111;
        10'd299   : cube_lut_0  = 14'b01101010111111;
        10'd300   : cube_lut_0  = 14'b01101011000110;
        10'd301   : cube_lut_0  = 14'b01101011001110;
        10'd302   : cube_lut_0  = 14'b01101011010110;
        10'd303   : cube_lut_0  = 14'b01101011011101;
        10'd304   : cube_lut_0  = 14'b01101011100101;
        10'd305   : cube_lut_0  = 14'b01101011101100;
        10'd306   : cube_lut_0  = 14'b01101011110100;
        10'd307   : cube_lut_0  = 14'b01101011111011;
        10'd308   : cube_lut_0  = 14'b01101100000011;
        10'd309   : cube_lut_0  = 14'b01101100001010;
        10'd310   : cube_lut_0  = 14'b01101100010010;
        10'd311   : cube_lut_0  = 14'b01101100011001;
        10'd312   : cube_lut_0  = 14'b01101100100001;
        10'd313   : cube_lut_0  = 14'b01101100101000;
        10'd314   : cube_lut_0  = 14'b01101100110000;
        10'd315   : cube_lut_0  = 14'b01101100110111;
        10'd316   : cube_lut_0  = 14'b01101100111110;
        10'd317   : cube_lut_0  = 14'b01101101000110;
        10'd318   : cube_lut_0  = 14'b01101101001101;
        10'd319   : cube_lut_0  = 14'b01101101010100;
        10'd320   : cube_lut_0  = 14'b01101101011100;
        10'd321   : cube_lut_0  = 14'b01101101100011;
        10'd322   : cube_lut_0  = 14'b01101101101010;
        10'd323   : cube_lut_0  = 14'b01101101110001;
        10'd324   : cube_lut_0  = 14'b01101101111001;
        10'd325   : cube_lut_0  = 14'b01101110000000;
        10'd326   : cube_lut_0  = 14'b01101110000111;
        10'd327   : cube_lut_0  = 14'b01101110001110;
        10'd328   : cube_lut_0  = 14'b01101110010101;
        10'd329   : cube_lut_0  = 14'b01101110011101;
        10'd330   : cube_lut_0  = 14'b01101110100100;
        10'd331   : cube_lut_0  = 14'b01101110101011;
        10'd332   : cube_lut_0  = 14'b01101110110010;
        10'd333   : cube_lut_0  = 14'b01101110111001;
        10'd334   : cube_lut_0  = 14'b01101111000000;
        10'd335   : cube_lut_0  = 14'b01101111000111;
        10'd336   : cube_lut_0  = 14'b01101111001110;
        10'd337   : cube_lut_0  = 14'b01101111010101;
        10'd338   : cube_lut_0  = 14'b01101111011100;
        10'd339   : cube_lut_0  = 14'b01101111100100;
        10'd340   : cube_lut_0  = 14'b01101111101011;
        10'd341   : cube_lut_0  = 14'b01101111110010;
        10'd342   : cube_lut_0  = 14'b01101111111001;
        10'd343   : cube_lut_0  = 14'b01110000000000;
        10'd344   : cube_lut_0  = 14'b01110000000110;
        10'd345   : cube_lut_0  = 14'b01110000001101;
        10'd346   : cube_lut_0  = 14'b01110000010100;
        10'd347   : cube_lut_0  = 14'b01110000011011;
        10'd348   : cube_lut_0  = 14'b01110000100010;
        10'd349   : cube_lut_0  = 14'b01110000101001;
        10'd350   : cube_lut_0  = 14'b01110000110000;
        10'd351   : cube_lut_0  = 14'b01110000110111;
        10'd352   : cube_lut_0  = 14'b01110000111110;
        10'd353   : cube_lut_0  = 14'b01110001000100;
        10'd354   : cube_lut_0  = 14'b01110001001011;
        10'd355   : cube_lut_0  = 14'b01110001010010;
        10'd356   : cube_lut_0  = 14'b01110001011001;
        10'd357   : cube_lut_0  = 14'b01110001100000;
        10'd358   : cube_lut_0  = 14'b01110001100111;
        10'd359   : cube_lut_0  = 14'b01110001101101;
        10'd360   : cube_lut_0  = 14'b01110001110100;
        10'd361   : cube_lut_0  = 14'b01110001111011;
        10'd362   : cube_lut_0  = 14'b01110010000001;
        10'd363   : cube_lut_0  = 14'b01110010001000;
        10'd364   : cube_lut_0  = 14'b01110010001111;
        10'd365   : cube_lut_0  = 14'b01110010010110;
        10'd366   : cube_lut_0  = 14'b01110010011100;
        10'd367   : cube_lut_0  = 14'b01110010100011;
        10'd368   : cube_lut_0  = 14'b01110010101010;
        10'd369   : cube_lut_0  = 14'b01110010110000;
        10'd370   : cube_lut_0  = 14'b01110010110111;
        10'd371   : cube_lut_0  = 14'b01110010111101;
        10'd372   : cube_lut_0  = 14'b01110011000100;
        10'd373   : cube_lut_0  = 14'b01110011001011;
        10'd374   : cube_lut_0  = 14'b01110011010001;
        10'd375   : cube_lut_0  = 14'b01110011011000;
        10'd376   : cube_lut_0  = 14'b01110011011110;
        10'd377   : cube_lut_0  = 14'b01110011100101;
        10'd378   : cube_lut_0  = 14'b01110011101011;
        10'd379   : cube_lut_0  = 14'b01110011110010;
        10'd380   : cube_lut_0  = 14'b01110011111000;
        10'd381   : cube_lut_0  = 14'b01110011111111;
        10'd382   : cube_lut_0  = 14'b01110100000101;
        10'd383   : cube_lut_0  = 14'b01110100001100;
        10'd384   : cube_lut_0  = 14'b01110100010010;
        10'd385   : cube_lut_0  = 14'b01110100011001;
        10'd386   : cube_lut_0  = 14'b01110100011111;
        10'd387   : cube_lut_0  = 14'b01110100100110;
        10'd388   : cube_lut_0  = 14'b01110100101100;
        10'd389   : cube_lut_0  = 14'b01110100110011;
        10'd390   : cube_lut_0  = 14'b01110100111001;
        10'd391   : cube_lut_0  = 14'b01110100111111;
        10'd392   : cube_lut_0  = 14'b01110101000110;
        10'd393   : cube_lut_0  = 14'b01110101001100;
        10'd394   : cube_lut_0  = 14'b01110101010010;
        10'd395   : cube_lut_0  = 14'b01110101011001;
        10'd396   : cube_lut_0  = 14'b01110101011111;
        10'd397   : cube_lut_0  = 14'b01110101100101;
        10'd398   : cube_lut_0  = 14'b01110101101100;
        10'd399   : cube_lut_0  = 14'b01110101110010;
        10'd400   : cube_lut_0  = 14'b01110101111000;
        10'd401   : cube_lut_0  = 14'b01110101111111;
        10'd402   : cube_lut_0  = 14'b01110110000101;
        10'd403   : cube_lut_0  = 14'b01110110001011;
        10'd404   : cube_lut_0  = 14'b01110110010001;
        10'd405   : cube_lut_0  = 14'b01110110011000;
        10'd406   : cube_lut_0  = 14'b01110110011110;
        10'd407   : cube_lut_0  = 14'b01110110100100;
        10'd408   : cube_lut_0  = 14'b01110110101010;
        10'd409   : cube_lut_0  = 14'b01110110110001;
        10'd410   : cube_lut_0  = 14'b01110110110111;
        10'd411   : cube_lut_0  = 14'b01110110111101;
        10'd412   : cube_lut_0  = 14'b01110111000011;
        10'd413   : cube_lut_0  = 14'b01110111001001;
        10'd414   : cube_lut_0  = 14'b01110111001111;
        10'd415   : cube_lut_0  = 14'b01110111010110;
        10'd416   : cube_lut_0  = 14'b01110111011100;
        10'd417   : cube_lut_0  = 14'b01110111100010;
        10'd418   : cube_lut_0  = 14'b01110111101000;
        10'd419   : cube_lut_0  = 14'b01110111101110;
        10'd420   : cube_lut_0  = 14'b01110111110100;
        10'd421   : cube_lut_0  = 14'b01110111111010;
        10'd422   : cube_lut_0  = 14'b01111000000000;
        10'd423   : cube_lut_0  = 14'b01111000000110;
        10'd424   : cube_lut_0  = 14'b01111000001100;
        10'd425   : cube_lut_0  = 14'b01111000010010;
        10'd426   : cube_lut_0  = 14'b01111000011000;
        10'd427   : cube_lut_0  = 14'b01111000011110;
        10'd428   : cube_lut_0  = 14'b01111000100100;
        10'd429   : cube_lut_0  = 14'b01111000101010;
        10'd430   : cube_lut_0  = 14'b01111000110000;
        10'd431   : cube_lut_0  = 14'b01111000110110;
        10'd432   : cube_lut_0  = 14'b01111000111100;
        10'd433   : cube_lut_0  = 14'b01111001000010;
        10'd434   : cube_lut_0  = 14'b01111001001000;
        10'd435   : cube_lut_0  = 14'b01111001001110;
        10'd436   : cube_lut_0  = 14'b01111001010100;
        10'd437   : cube_lut_0  = 14'b01111001011010;
        10'd438   : cube_lut_0  = 14'b01111001100000;
        10'd439   : cube_lut_0  = 14'b01111001100110;
        10'd440   : cube_lut_0  = 14'b01111001101100;
        10'd441   : cube_lut_0  = 14'b01111001110010;
        10'd442   : cube_lut_0  = 14'b01111001111000;
        10'd443   : cube_lut_0  = 14'b01111001111110;
        10'd444   : cube_lut_0  = 14'b01111010000011;
        10'd445   : cube_lut_0  = 14'b01111010001001;
        10'd446   : cube_lut_0  = 14'b01111010001111;
        10'd447   : cube_lut_0  = 14'b01111010010101;
        10'd448   : cube_lut_0  = 14'b01111010011011;
        10'd449   : cube_lut_0  = 14'b01111010100001;
        10'd450   : cube_lut_0  = 14'b01111010100111;
        10'd451   : cube_lut_0  = 14'b01111010101100;
        10'd452   : cube_lut_0  = 14'b01111010110010;
        10'd453   : cube_lut_0  = 14'b01111010111000;
        10'd454   : cube_lut_0  = 14'b01111010111110;
        10'd455   : cube_lut_0  = 14'b01111011000011;
        10'd456   : cube_lut_0  = 14'b01111011001001;
        10'd457   : cube_lut_0  = 14'b01111011001111;
        10'd458   : cube_lut_0  = 14'b01111011010101;
        10'd459   : cube_lut_0  = 14'b01111011011010;
        10'd460   : cube_lut_0  = 14'b01111011100000;
        10'd461   : cube_lut_0  = 14'b01111011100110;
        10'd462   : cube_lut_0  = 14'b01111011101100;
        10'd463   : cube_lut_0  = 14'b01111011110001;
        10'd464   : cube_lut_0  = 14'b01111011110111;
        10'd465   : cube_lut_0  = 14'b01111011111101;
        10'd466   : cube_lut_0  = 14'b01111100000010;
        10'd467   : cube_lut_0  = 14'b01111100001000;
        10'd468   : cube_lut_0  = 14'b01111100001110;
        10'd469   : cube_lut_0  = 14'b01111100010011;
        10'd470   : cube_lut_0  = 14'b01111100011001;
        10'd471   : cube_lut_0  = 14'b01111100011111;
        10'd472   : cube_lut_0  = 14'b01111100100100;
        10'd473   : cube_lut_0  = 14'b01111100101010;
        10'd474   : cube_lut_0  = 14'b01111100110000;
        10'd475   : cube_lut_0  = 14'b01111100110101;
        10'd476   : cube_lut_0  = 14'b01111100111011;
        10'd477   : cube_lut_0  = 14'b01111101000000;
        10'd478   : cube_lut_0  = 14'b01111101000110;
        10'd479   : cube_lut_0  = 14'b01111101001100;
        10'd480   : cube_lut_0  = 14'b01111101010001;
        10'd481   : cube_lut_0  = 14'b01111101010111;
        10'd482   : cube_lut_0  = 14'b01111101011100;
        10'd483   : cube_lut_0  = 14'b01111101100010;
        10'd484   : cube_lut_0  = 14'b01111101100111;
        10'd485   : cube_lut_0  = 14'b01111101101101;
        10'd486   : cube_lut_0  = 14'b01111101110010;
        10'd487   : cube_lut_0  = 14'b01111101111000;
        10'd488   : cube_lut_0  = 14'b01111101111101;
        10'd489   : cube_lut_0  = 14'b01111110000011;
        10'd490   : cube_lut_0  = 14'b01111110001000;
        10'd491   : cube_lut_0  = 14'b01111110001110;
        10'd492   : cube_lut_0  = 14'b01111110010011;
        10'd493   : cube_lut_0  = 14'b01111110011001;
        10'd494   : cube_lut_0  = 14'b01111110011110;
        10'd495   : cube_lut_0  = 14'b01111110100100;
        10'd496   : cube_lut_0  = 14'b01111110101001;
        10'd497   : cube_lut_0  = 14'b01111110101111;
        10'd498   : cube_lut_0  = 14'b01111110110100;
        10'd499   : cube_lut_0  = 14'b01111110111010;
        10'd500   : cube_lut_0  = 14'b01111110111111;
        10'd501   : cube_lut_0  = 14'b01111111000100;
        10'd502   : cube_lut_0  = 14'b01111111001010;
        10'd503   : cube_lut_0  = 14'b01111111001111;
        10'd504   : cube_lut_0  = 14'b01111111010101;
        10'd505   : cube_lut_0  = 14'b01111111011010;
        10'd506   : cube_lut_0  = 14'b01111111011111;
        10'd507   : cube_lut_0  = 14'b01111111100101;
        10'd508   : cube_lut_0  = 14'b01111111101010;
        10'd509   : cube_lut_0  = 14'b01111111101111;
        10'd510   : cube_lut_0  = 14'b01111111110101;
        10'd511   : cube_lut_0  = 14'b01111111111010;
        10'd512   : cube_lut_0  = 14'b10000000000000;
        10'd513   : cube_lut_0  = 14'b10000000000101;
        10'd514   : cube_lut_0  = 14'b10000000001010;
        10'd515   : cube_lut_0  = 14'b10000000001111;
        10'd516   : cube_lut_0  = 14'b10000000010101;
        10'd517   : cube_lut_0  = 14'b10000000011010;
        10'd518   : cube_lut_0  = 14'b10000000011111;
        10'd519   : cube_lut_0  = 14'b10000000100101;
        10'd520   : cube_lut_0  = 14'b10000000101010;
        10'd521   : cube_lut_0  = 14'b10000000101111;
        10'd522   : cube_lut_0  = 14'b10000000110100;
        10'd523   : cube_lut_0  = 14'b10000000111010;
        10'd524   : cube_lut_0  = 14'b10000000111111;
        10'd525   : cube_lut_0  = 14'b10000001000100;
        10'd526   : cube_lut_0  = 14'b10000001001001;
        10'd527   : cube_lut_0  = 14'b10000001001111;
        10'd528   : cube_lut_0  = 14'b10000001010100;
        10'd529   : cube_lut_0  = 14'b10000001011001;
        10'd530   : cube_lut_0  = 14'b10000001011110;
        10'd531   : cube_lut_0  = 14'b10000001100100;
        10'd532   : cube_lut_0  = 14'b10000001101001;
        10'd533   : cube_lut_0  = 14'b10000001101110;
        10'd534   : cube_lut_0  = 14'b10000001110011;
        10'd535   : cube_lut_0  = 14'b10000001111000;
        10'd536   : cube_lut_0  = 14'b10000001111110;
        10'd537   : cube_lut_0  = 14'b10000010000011;
        10'd538   : cube_lut_0  = 14'b10000010001000;
        10'd539   : cube_lut_0  = 14'b10000010001101;
        10'd540   : cube_lut_0  = 14'b10000010010010;
        10'd541   : cube_lut_0  = 14'b10000010010111;
        10'd542   : cube_lut_0  = 14'b10000010011100;
        10'd543   : cube_lut_0  = 14'b10000010100010;
        10'd544   : cube_lut_0  = 14'b10000010100111;
        10'd545   : cube_lut_0  = 14'b10000010101100;
        10'd546   : cube_lut_0  = 14'b10000010110001;
        10'd547   : cube_lut_0  = 14'b10000010110110;
        10'd548   : cube_lut_0  = 14'b10000010111011;
        10'd549   : cube_lut_0  = 14'b10000011000000;
        10'd550   : cube_lut_0  = 14'b10000011000101;
        10'd551   : cube_lut_0  = 14'b10000011001010;
        10'd552   : cube_lut_0  = 14'b10000011010000;
        10'd553   : cube_lut_0  = 14'b10000011010101;
        10'd554   : cube_lut_0  = 14'b10000011011010;
        10'd555   : cube_lut_0  = 14'b10000011011111;
        10'd556   : cube_lut_0  = 14'b10000011100100;
        10'd557   : cube_lut_0  = 14'b10000011101001;
        10'd558   : cube_lut_0  = 14'b10000011101110;
        10'd559   : cube_lut_0  = 14'b10000011110011;
        10'd560   : cube_lut_0  = 14'b10000011111000;
        10'd561   : cube_lut_0  = 14'b10000011111101;
        10'd562   : cube_lut_0  = 14'b10000100000010;
        10'd563   : cube_lut_0  = 14'b10000100000111;
        10'd564   : cube_lut_0  = 14'b10000100001100;
        10'd565   : cube_lut_0  = 14'b10000100010001;
        10'd566   : cube_lut_0  = 14'b10000100010110;
        10'd567   : cube_lut_0  = 14'b10000100011011;
        10'd568   : cube_lut_0  = 14'b10000100100000;
        10'd569   : cube_lut_0  = 14'b10000100100101;
        10'd570   : cube_lut_0  = 14'b10000100101010;
        10'd571   : cube_lut_0  = 14'b10000100101111;
        10'd572   : cube_lut_0  = 14'b10000100110100;
        10'd573   : cube_lut_0  = 14'b10000100111001;
        10'd574   : cube_lut_0  = 14'b10000100111110;
        10'd575   : cube_lut_0  = 14'b10000101000011;
        10'd576   : cube_lut_0  = 14'b10000101001000;
        10'd577   : cube_lut_0  = 14'b10000101001100;
        10'd578   : cube_lut_0  = 14'b10000101010001;
        10'd579   : cube_lut_0  = 14'b10000101010110;
        10'd580   : cube_lut_0  = 14'b10000101011011;
        10'd581   : cube_lut_0  = 14'b10000101100000;
        10'd582   : cube_lut_0  = 14'b10000101100101;
        10'd583   : cube_lut_0  = 14'b10000101101010;
        10'd584   : cube_lut_0  = 14'b10000101101111;
        10'd585   : cube_lut_0  = 14'b10000101110100;
        10'd586   : cube_lut_0  = 14'b10000101111001;
        10'd587   : cube_lut_0  = 14'b10000101111101;
        10'd588   : cube_lut_0  = 14'b10000110000010;
        10'd589   : cube_lut_0  = 14'b10000110000111;
        10'd590   : cube_lut_0  = 14'b10000110001100;
        10'd591   : cube_lut_0  = 14'b10000110010001;
        10'd592   : cube_lut_0  = 14'b10000110010110;
        10'd593   : cube_lut_0  = 14'b10000110011011;
        10'd594   : cube_lut_0  = 14'b10000110011111;
        10'd595   : cube_lut_0  = 14'b10000110100100;
        10'd596   : cube_lut_0  = 14'b10000110101001;
        10'd597   : cube_lut_0  = 14'b10000110101110;
        10'd598   : cube_lut_0  = 14'b10000110110011;
        10'd599   : cube_lut_0  = 14'b10000110110111;
        10'd600   : cube_lut_0  = 14'b10000110111100;
        10'd601   : cube_lut_0  = 14'b10000111000001;
        10'd602   : cube_lut_0  = 14'b10000111000110;
        10'd603   : cube_lut_0  = 14'b10000111001011;
        10'd604   : cube_lut_0  = 14'b10000111001111;
        10'd605   : cube_lut_0  = 14'b10000111010100;
        10'd606   : cube_lut_0  = 14'b10000111011001;
        10'd607   : cube_lut_0  = 14'b10000111011110;
        10'd608   : cube_lut_0  = 14'b10000111100010;
        10'd609   : cube_lut_0  = 14'b10000111100111;
        10'd610   : cube_lut_0  = 14'b10000111101100;
        10'd611   : cube_lut_0  = 14'b10000111110001;
        10'd612   : cube_lut_0  = 14'b10000111110101;
        10'd613   : cube_lut_0  = 14'b10000111111010;
        10'd614   : cube_lut_0  = 14'b10000111111111;
        10'd615   : cube_lut_0  = 14'b10001000000100;
        10'd616   : cube_lut_0  = 14'b10001000001000;
        10'd617   : cube_lut_0  = 14'b10001000001101;
        10'd618   : cube_lut_0  = 14'b10001000010010;
        10'd619   : cube_lut_0  = 14'b10001000010110;
        10'd620   : cube_lut_0  = 14'b10001000011011;
        10'd621   : cube_lut_0  = 14'b10001000100000;
        10'd622   : cube_lut_0  = 14'b10001000100101;
        10'd623   : cube_lut_0  = 14'b10001000101001;
        10'd624   : cube_lut_0  = 14'b10001000101110;
        10'd625   : cube_lut_0  = 14'b10001000110011;
        10'd626   : cube_lut_0  = 14'b10001000110111;
        10'd627   : cube_lut_0  = 14'b10001000111100;
        10'd628   : cube_lut_0  = 14'b10001001000001;
        10'd629   : cube_lut_0  = 14'b10001001000101;
        10'd630   : cube_lut_0  = 14'b10001001001010;
        10'd631   : cube_lut_0  = 14'b10001001001111;
        10'd632   : cube_lut_0  = 14'b10001001010011;
        10'd633   : cube_lut_0  = 14'b10001001011000;
        10'd634   : cube_lut_0  = 14'b10001001011100;
        10'd635   : cube_lut_0  = 14'b10001001100001;
        10'd636   : cube_lut_0  = 14'b10001001100110;
        10'd637   : cube_lut_0  = 14'b10001001101010;
        10'd638   : cube_lut_0  = 14'b10001001101111;
        10'd639   : cube_lut_0  = 14'b10001001110011;
        10'd640   : cube_lut_0  = 14'b10001001111000;
        10'd641   : cube_lut_0  = 14'b10001001111101;
        10'd642   : cube_lut_0  = 14'b10001010000001;
        10'd643   : cube_lut_0  = 14'b10001010000110;
        10'd644   : cube_lut_0  = 14'b10001010001010;
        10'd645   : cube_lut_0  = 14'b10001010001111;
        10'd646   : cube_lut_0  = 14'b10001010010100;
        10'd647   : cube_lut_0  = 14'b10001010011000;
        10'd648   : cube_lut_0  = 14'b10001010011101;
        10'd649   : cube_lut_0  = 14'b10001010100001;
        10'd650   : cube_lut_0  = 14'b10001010100110;
        10'd651   : cube_lut_0  = 14'b10001010101010;
        10'd652   : cube_lut_0  = 14'b10001010101111;
        10'd653   : cube_lut_0  = 14'b10001010110011;
        10'd654   : cube_lut_0  = 14'b10001010111000;
        10'd655   : cube_lut_0  = 14'b10001010111100;
        10'd656   : cube_lut_0  = 14'b10001011000001;
        10'd657   : cube_lut_0  = 14'b10001011000110;
        10'd658   : cube_lut_0  = 14'b10001011001010;
        10'd659   : cube_lut_0  = 14'b10001011001111;
        10'd660   : cube_lut_0  = 14'b10001011010011;
        10'd661   : cube_lut_0  = 14'b10001011011000;
        10'd662   : cube_lut_0  = 14'b10001011011100;
        10'd663   : cube_lut_0  = 14'b10001011100001;
        10'd664   : cube_lut_0  = 14'b10001011100101;
        10'd665   : cube_lut_0  = 14'b10001011101010;
        10'd666   : cube_lut_0  = 14'b10001011101110;
        10'd667   : cube_lut_0  = 14'b10001011110010;
        10'd668   : cube_lut_0  = 14'b10001011110111;
        10'd669   : cube_lut_0  = 14'b10001011111011;
        10'd670   : cube_lut_0  = 14'b10001100000000;
        10'd671   : cube_lut_0  = 14'b10001100000100;
        10'd672   : cube_lut_0  = 14'b10001100001001;
        10'd673   : cube_lut_0  = 14'b10001100001101;
        10'd674   : cube_lut_0  = 14'b10001100010010;
        10'd675   : cube_lut_0  = 14'b10001100010110;
        10'd676   : cube_lut_0  = 14'b10001100011011;
        10'd677   : cube_lut_0  = 14'b10001100011111;
        10'd678   : cube_lut_0  = 14'b10001100100011;
        10'd679   : cube_lut_0  = 14'b10001100101000;
        10'd680   : cube_lut_0  = 14'b10001100101100;
        10'd681   : cube_lut_0  = 14'b10001100110001;
        10'd682   : cube_lut_0  = 14'b10001100110101;
        10'd683   : cube_lut_0  = 14'b10001100111001;
        10'd684   : cube_lut_0  = 14'b10001100111110;
        10'd685   : cube_lut_0  = 14'b10001101000010;
        10'd686   : cube_lut_0  = 14'b10001101000111;
        10'd687   : cube_lut_0  = 14'b10001101001011;
        10'd688   : cube_lut_0  = 14'b10001101001111;
        10'd689   : cube_lut_0  = 14'b10001101010100;
        10'd690   : cube_lut_0  = 14'b10001101011000;
        10'd691   : cube_lut_0  = 14'b10001101011101;
        10'd692   : cube_lut_0  = 14'b10001101100001;
        10'd693   : cube_lut_0  = 14'b10001101100101;
        10'd694   : cube_lut_0  = 14'b10001101101010;
        10'd695   : cube_lut_0  = 14'b10001101101110;
        10'd696   : cube_lut_0  = 14'b10001101110010;
        10'd697   : cube_lut_0  = 14'b10001101110111;
        10'd698   : cube_lut_0  = 14'b10001101111011;
        10'd699   : cube_lut_0  = 14'b10001101111111;
        10'd700   : cube_lut_0  = 14'b10001110000100;
        10'd701   : cube_lut_0  = 14'b10001110001000;
        10'd702   : cube_lut_0  = 14'b10001110001100;
        10'd703   : cube_lut_0  = 14'b10001110010001;
        10'd704   : cube_lut_0  = 14'b10001110010101;
        10'd705   : cube_lut_0  = 14'b10001110011001;
        10'd706   : cube_lut_0  = 14'b10001110011110;
        10'd707   : cube_lut_0  = 14'b10001110100010;
        10'd708   : cube_lut_0  = 14'b10001110100110;
        10'd709   : cube_lut_0  = 14'b10001110101010;
        10'd710   : cube_lut_0  = 14'b10001110101111;
        10'd711   : cube_lut_0  = 14'b10001110110011;
        10'd712   : cube_lut_0  = 14'b10001110110111;
        10'd713   : cube_lut_0  = 14'b10001110111100;
        10'd714   : cube_lut_0  = 14'b10001111000000;
        10'd715   : cube_lut_0  = 14'b10001111000100;
        10'd716   : cube_lut_0  = 14'b10001111001000;
        10'd717   : cube_lut_0  = 14'b10001111001101;
        10'd718   : cube_lut_0  = 14'b10001111010001;
        10'd719   : cube_lut_0  = 14'b10001111010101;
        10'd720   : cube_lut_0  = 14'b10001111011001;
        10'd721   : cube_lut_0  = 14'b10001111011110;
        10'd722   : cube_lut_0  = 14'b10001111100010;
        10'd723   : cube_lut_0  = 14'b10001111100110;
        10'd724   : cube_lut_0  = 14'b10001111101010;
        10'd725   : cube_lut_0  = 14'b10001111101111;
        10'd726   : cube_lut_0  = 14'b10001111110011;
        10'd727   : cube_lut_0  = 14'b10001111110111;
        10'd728   : cube_lut_0  = 14'b10001111111011;
        10'd729   : cube_lut_0  = 14'b10010000000000;
        10'd730   : cube_lut_0  = 14'b10010000000100;
        10'd731   : cube_lut_0  = 14'b10010000001000;
        10'd732   : cube_lut_0  = 14'b10010000001100;
        10'd733   : cube_lut_0  = 14'b10010000010000;
        10'd734   : cube_lut_0  = 14'b10010000010101;
        10'd735   : cube_lut_0  = 14'b10010000011001;
        10'd736   : cube_lut_0  = 14'b10010000011101;
        10'd737   : cube_lut_0  = 14'b10010000100001;
        10'd738   : cube_lut_0  = 14'b10010000100101;
        10'd739   : cube_lut_0  = 14'b10010000101001;
        10'd740   : cube_lut_0  = 14'b10010000101110;
        10'd741   : cube_lut_0  = 14'b10010000110010;
        10'd742   : cube_lut_0  = 14'b10010000110110;
        10'd743   : cube_lut_0  = 14'b10010000111010;
        10'd744   : cube_lut_0  = 14'b10010000111110;
        10'd745   : cube_lut_0  = 14'b10010001000010;
        10'd746   : cube_lut_0  = 14'b10010001000111;
        10'd747   : cube_lut_0  = 14'b10010001001011;
        10'd748   : cube_lut_0  = 14'b10010001001111;
        10'd749   : cube_lut_0  = 14'b10010001010011;
        10'd750   : cube_lut_0  = 14'b10010001010111;
        10'd751   : cube_lut_0  = 14'b10010001011011;
        10'd752   : cube_lut_0  = 14'b10010001011111;
        10'd753   : cube_lut_0  = 14'b10010001100100;
        10'd754   : cube_lut_0  = 14'b10010001101000;
        10'd755   : cube_lut_0  = 14'b10010001101100;
        10'd756   : cube_lut_0  = 14'b10010001110000;
        10'd757   : cube_lut_0  = 14'b10010001110100;
        10'd758   : cube_lut_0  = 14'b10010001111000;
        10'd759   : cube_lut_0  = 14'b10010001111100;
        10'd760   : cube_lut_0  = 14'b10010010000000;
        10'd761   : cube_lut_0  = 14'b10010010000100;
        10'd762   : cube_lut_0  = 14'b10010010001001;
        10'd763   : cube_lut_0  = 14'b10010010001101;
        10'd764   : cube_lut_0  = 14'b10010010010001;
        10'd765   : cube_lut_0  = 14'b10010010010101;
        10'd766   : cube_lut_0  = 14'b10010010011001;
        10'd767   : cube_lut_0  = 14'b10010010011101;
        10'd768   : cube_lut_0  = 14'b10010010100001;
        10'd769   : cube_lut_0  = 14'b10010010100101;
        10'd770   : cube_lut_0  = 14'b10010010101001;
        10'd771   : cube_lut_0  = 14'b10010010101101;
        10'd772   : cube_lut_0  = 14'b10010010110001;
        10'd773   : cube_lut_0  = 14'b10010010110101;
        10'd774   : cube_lut_0  = 14'b10010010111001;
        10'd775   : cube_lut_0  = 14'b10010010111101;
        10'd776   : cube_lut_0  = 14'b10010011000001;
        10'd777   : cube_lut_0  = 14'b10010011000101;
        10'd778   : cube_lut_0  = 14'b10010011001010;
        10'd779   : cube_lut_0  = 14'b10010011001110;
        10'd780   : cube_lut_0  = 14'b10010011010010;
        10'd781   : cube_lut_0  = 14'b10010011010110;
        10'd782   : cube_lut_0  = 14'b10010011011010;
        10'd783   : cube_lut_0  = 14'b10010011011110;
        10'd784   : cube_lut_0  = 14'b10010011100010;
        10'd785   : cube_lut_0  = 14'b10010011100110;
        10'd786   : cube_lut_0  = 14'b10010011101010;
        10'd787   : cube_lut_0  = 14'b10010011101110;
        10'd788   : cube_lut_0  = 14'b10010011110010;
        10'd789   : cube_lut_0  = 14'b10010011110110;
        10'd790   : cube_lut_0  = 14'b10010011111010;
        10'd791   : cube_lut_0  = 14'b10010011111110;
        10'd792   : cube_lut_0  = 14'b10010100000010;
        10'd793   : cube_lut_0  = 14'b10010100000110;
        10'd794   : cube_lut_0  = 14'b10010100001010;
        10'd795   : cube_lut_0  = 14'b10010100001110;
        10'd796   : cube_lut_0  = 14'b10010100010010;
        10'd797   : cube_lut_0  = 14'b10010100010110;
        10'd798   : cube_lut_0  = 14'b10010100011010;
        10'd799   : cube_lut_0  = 14'b10010100011110;
        10'd800   : cube_lut_0  = 14'b10010100100001;
        10'd801   : cube_lut_0  = 14'b10010100100101;
        10'd802   : cube_lut_0  = 14'b10010100101001;
        10'd803   : cube_lut_0  = 14'b10010100101101;
        10'd804   : cube_lut_0  = 14'b10010100110001;
        10'd805   : cube_lut_0  = 14'b10010100110101;
        10'd806   : cube_lut_0  = 14'b10010100111001;
        10'd807   : cube_lut_0  = 14'b10010100111101;
        10'd808   : cube_lut_0  = 14'b10010101000001;
        10'd809   : cube_lut_0  = 14'b10010101000101;
        10'd810   : cube_lut_0  = 14'b10010101001001;
        10'd811   : cube_lut_0  = 14'b10010101001101;
        10'd812   : cube_lut_0  = 14'b10010101010001;
        10'd813   : cube_lut_0  = 14'b10010101010101;
        10'd814   : cube_lut_0  = 14'b10010101011001;
        10'd815   : cube_lut_0  = 14'b10010101011101;
        10'd816   : cube_lut_0  = 14'b10010101100000;
        10'd817   : cube_lut_0  = 14'b10010101100100;
        10'd818   : cube_lut_0  = 14'b10010101101000;
        10'd819   : cube_lut_0  = 14'b10010101101100;
        10'd820   : cube_lut_0  = 14'b10010101110000;
        10'd821   : cube_lut_0  = 14'b10010101110100;
        10'd822   : cube_lut_0  = 14'b10010101111000;
        10'd823   : cube_lut_0  = 14'b10010101111100;
        10'd824   : cube_lut_0  = 14'b10010110000000;
        10'd825   : cube_lut_0  = 14'b10010110000011;
        10'd826   : cube_lut_0  = 14'b10010110000111;
        10'd827   : cube_lut_0  = 14'b10010110001011;
        10'd828   : cube_lut_0  = 14'b10010110001111;
        10'd829   : cube_lut_0  = 14'b10010110010011;
        10'd830   : cube_lut_0  = 14'b10010110010111;
        10'd831   : cube_lut_0  = 14'b10010110011011;
        10'd832   : cube_lut_0  = 14'b10010110011111;
        10'd833   : cube_lut_0  = 14'b10010110100010;
        10'd834   : cube_lut_0  = 14'b10010110100110;
        10'd835   : cube_lut_0  = 14'b10010110101010;
        10'd836   : cube_lut_0  = 14'b10010110101110;
        10'd837   : cube_lut_0  = 14'b10010110110010;
        10'd838   : cube_lut_0  = 14'b10010110110110;
        10'd839   : cube_lut_0  = 14'b10010110111010;
        10'd840   : cube_lut_0  = 14'b10010110111101;
        10'd841   : cube_lut_0  = 14'b10010111000001;
        10'd842   : cube_lut_0  = 14'b10010111000101;
        10'd843   : cube_lut_0  = 14'b10010111001001;
        10'd844   : cube_lut_0  = 14'b10010111001101;
        10'd845   : cube_lut_0  = 14'b10010111010000;
        10'd846   : cube_lut_0  = 14'b10010111010100;
        10'd847   : cube_lut_0  = 14'b10010111011000;
        10'd848   : cube_lut_0  = 14'b10010111011100;
        10'd849   : cube_lut_0  = 14'b10010111100000;
        10'd850   : cube_lut_0  = 14'b10010111100100;
        10'd851   : cube_lut_0  = 14'b10010111100111;
        10'd852   : cube_lut_0  = 14'b10010111101011;
        10'd853   : cube_lut_0  = 14'b10010111101111;
        10'd854   : cube_lut_0  = 14'b10010111110011;
        10'd855   : cube_lut_0  = 14'b10010111110111;
        10'd856   : cube_lut_0  = 14'b10010111111010;
        10'd857   : cube_lut_0  = 14'b10010111111110;
        10'd858   : cube_lut_0  = 14'b10011000000010;
        10'd859   : cube_lut_0  = 14'b10011000000110;
        10'd860   : cube_lut_0  = 14'b10011000001001;
        10'd861   : cube_lut_0  = 14'b10011000001101;
        10'd862   : cube_lut_0  = 14'b10011000010001;
        10'd863   : cube_lut_0  = 14'b10011000010101;
        10'd864   : cube_lut_0  = 14'b10011000011000;
        10'd865   : cube_lut_0  = 14'b10011000011100;
        10'd866   : cube_lut_0  = 14'b10011000100000;
        10'd867   : cube_lut_0  = 14'b10011000100100;
        10'd868   : cube_lut_0  = 14'b10011000101000;
        10'd869   : cube_lut_0  = 14'b10011000101011;
        10'd870   : cube_lut_0  = 14'b10011000101111;
        10'd871   : cube_lut_0  = 14'b10011000110011;
        10'd872   : cube_lut_0  = 14'b10011000110111;
        10'd873   : cube_lut_0  = 14'b10011000111010;
        10'd874   : cube_lut_0  = 14'b10011000111110;
        10'd875   : cube_lut_0  = 14'b10011001000010;
        10'd876   : cube_lut_0  = 14'b10011001000101;
        10'd877   : cube_lut_0  = 14'b10011001001001;
        10'd878   : cube_lut_0  = 14'b10011001001101;
        10'd879   : cube_lut_0  = 14'b10011001010001;
        10'd880   : cube_lut_0  = 14'b10011001010100;
        10'd881   : cube_lut_0  = 14'b10011001011000;
        10'd882   : cube_lut_0  = 14'b10011001011100;
        10'd883   : cube_lut_0  = 14'b10011001011111;
        10'd884   : cube_lut_0  = 14'b10011001100011;
        10'd885   : cube_lut_0  = 14'b10011001100111;
        10'd886   : cube_lut_0  = 14'b10011001101011;
        10'd887   : cube_lut_0  = 14'b10011001101110;
        10'd888   : cube_lut_0  = 14'b10011001110010;
        10'd889   : cube_lut_0  = 14'b10011001110110;
        10'd890   : cube_lut_0  = 14'b10011001111001;
        10'd891   : cube_lut_0  = 14'b10011001111101;
        10'd892   : cube_lut_0  = 14'b10011010000001;
        10'd893   : cube_lut_0  = 14'b10011010000100;
        10'd894   : cube_lut_0  = 14'b10011010001000;
        10'd895   : cube_lut_0  = 14'b10011010001100;
        10'd896   : cube_lut_0  = 14'b10011010001111;
        10'd897   : cube_lut_0  = 14'b10011010010011;
        10'd898   : cube_lut_0  = 14'b10011010010111;
        10'd899   : cube_lut_0  = 14'b10011010011010;
        10'd900   : cube_lut_0  = 14'b10011010011110;
        10'd901   : cube_lut_0  = 14'b10011010100010;
        10'd902   : cube_lut_0  = 14'b10011010100101;
        10'd903   : cube_lut_0  = 14'b10011010101001;
        10'd904   : cube_lut_0  = 14'b10011010101101;
        10'd905   : cube_lut_0  = 14'b10011010110000;
        10'd906   : cube_lut_0  = 14'b10011010110100;
        10'd907   : cube_lut_0  = 14'b10011010111000;
        10'd908   : cube_lut_0  = 14'b10011010111011;
        10'd909   : cube_lut_0  = 14'b10011010111111;
        10'd910   : cube_lut_0  = 14'b10011011000011;
        10'd911   : cube_lut_0  = 14'b10011011000110;
        10'd912   : cube_lut_0  = 14'b10011011001010;
        10'd913   : cube_lut_0  = 14'b10011011001101;
        10'd914   : cube_lut_0  = 14'b10011011010001;
        10'd915   : cube_lut_0  = 14'b10011011010101;
        10'd916   : cube_lut_0  = 14'b10011011011000;
        10'd917   : cube_lut_0  = 14'b10011011011100;
        10'd918   : cube_lut_0  = 14'b10011011100000;
        10'd919   : cube_lut_0  = 14'b10011011100011;
        10'd920   : cube_lut_0  = 14'b10011011100111;
        10'd921   : cube_lut_0  = 14'b10011011101010;
        10'd922   : cube_lut_0  = 14'b10011011101110;
        10'd923   : cube_lut_0  = 14'b10011011110010;
        10'd924   : cube_lut_0  = 14'b10011011110101;
        10'd925   : cube_lut_0  = 14'b10011011111001;
        10'd926   : cube_lut_0  = 14'b10011011111100;
        10'd927   : cube_lut_0  = 14'b10011100000000;
        10'd928   : cube_lut_0  = 14'b10011100000100;
        10'd929   : cube_lut_0  = 14'b10011100000111;
        10'd930   : cube_lut_0  = 14'b10011100001011;
        10'd931   : cube_lut_0  = 14'b10011100001110;
        10'd932   : cube_lut_0  = 14'b10011100010010;
        10'd933   : cube_lut_0  = 14'b10011100010110;
        10'd934   : cube_lut_0  = 14'b10011100011001;
        10'd935   : cube_lut_0  = 14'b10011100011101;
        10'd936   : cube_lut_0  = 14'b10011100100000;
        10'd937   : cube_lut_0  = 14'b10011100100100;
        10'd938   : cube_lut_0  = 14'b10011100100111;
        10'd939   : cube_lut_0  = 14'b10011100101011;
        10'd940   : cube_lut_0  = 14'b10011100101110;
        10'd941   : cube_lut_0  = 14'b10011100110010;
        10'd942   : cube_lut_0  = 14'b10011100110110;
        10'd943   : cube_lut_0  = 14'b10011100111001;
        10'd944   : cube_lut_0  = 14'b10011100111101;
        10'd945   : cube_lut_0  = 14'b10011101000000;
        10'd946   : cube_lut_0  = 14'b10011101000100;
        10'd947   : cube_lut_0  = 14'b10011101000111;
        10'd948   : cube_lut_0  = 14'b10011101001011;
        10'd949   : cube_lut_0  = 14'b10011101001110;
        10'd950   : cube_lut_0  = 14'b10011101010010;
        10'd951   : cube_lut_0  = 14'b10011101010101;
        10'd952   : cube_lut_0  = 14'b10011101011001;
        10'd953   : cube_lut_0  = 14'b10011101011100;
        10'd954   : cube_lut_0  = 14'b10011101100000;
        10'd955   : cube_lut_0  = 14'b10011101100100;
        10'd956   : cube_lut_0  = 14'b10011101100111;
        10'd957   : cube_lut_0  = 14'b10011101101011;
        10'd958   : cube_lut_0  = 14'b10011101101110;
        10'd959   : cube_lut_0  = 14'b10011101110010;
        10'd960   : cube_lut_0  = 14'b10011101110101;
        10'd961   : cube_lut_0  = 14'b10011101111001;
        10'd962   : cube_lut_0  = 14'b10011101111100;
        10'd963   : cube_lut_0  = 14'b10011110000000;
        10'd964   : cube_lut_0  = 14'b10011110000011;
        10'd965   : cube_lut_0  = 14'b10011110000111;
        10'd966   : cube_lut_0  = 14'b10011110001010;
        10'd967   : cube_lut_0  = 14'b10011110001110;
        10'd968   : cube_lut_0  = 14'b10011110010001;
        10'd969   : cube_lut_0  = 14'b10011110010101;
        10'd970   : cube_lut_0  = 14'b10011110011000;
        10'd971   : cube_lut_0  = 14'b10011110011100;
        10'd972   : cube_lut_0  = 14'b10011110011111;
        10'd973   : cube_lut_0  = 14'b10011110100010;
        10'd974   : cube_lut_0  = 14'b10011110100110;
        10'd975   : cube_lut_0  = 14'b10011110101001;
        10'd976   : cube_lut_0  = 14'b10011110101101;
        10'd977   : cube_lut_0  = 14'b10011110110000;
        10'd978   : cube_lut_0  = 14'b10011110110100;
        10'd979   : cube_lut_0  = 14'b10011110110111;
        10'd980   : cube_lut_0  = 14'b10011110111011;
        10'd981   : cube_lut_0  = 14'b10011110111110;
        10'd982   : cube_lut_0  = 14'b10011111000010;
        10'd983   : cube_lut_0  = 14'b10011111000101;
        10'd984   : cube_lut_0  = 14'b10011111001001;
        10'd985   : cube_lut_0  = 14'b10011111001100;
        10'd986   : cube_lut_0  = 14'b10011111001111;
        10'd987   : cube_lut_0  = 14'b10011111010011;
        10'd988   : cube_lut_0  = 14'b10011111010110;
        10'd989   : cube_lut_0  = 14'b10011111011010;
        10'd990   : cube_lut_0  = 14'b10011111011101;
        10'd991   : cube_lut_0  = 14'b10011111100001;
        10'd992   : cube_lut_0  = 14'b10011111100100;
        10'd993   : cube_lut_0  = 14'b10011111101000;
        10'd994   : cube_lut_0  = 14'b10011111101011;
        10'd995   : cube_lut_0  = 14'b10011111101110;
        10'd996   : cube_lut_0  = 14'b10011111110010;
        10'd997   : cube_lut_0  = 14'b10011111110101;
        10'd998   : cube_lut_0  = 14'b10011111111001;
        10'd999   : cube_lut_0  = 14'b10011111111100;
        10'd1000   : cube_lut_0 = 14'b10100000000000;
        10'd1001   : cube_lut_0 = 14'b10100000000011;
        10'd1002   : cube_lut_0 = 14'b10100000000110;
        10'd1003   : cube_lut_0 = 14'b10100000001010;
        10'd1004   : cube_lut_0 = 14'b10100000001101;
        10'd1005   : cube_lut_0 = 14'b10100000010001;
        10'd1006   : cube_lut_0 = 14'b10100000010100;
        10'd1007   : cube_lut_0 = 14'b10100000010111;
        10'd1008   : cube_lut_0 = 14'b10100000011011;
        10'd1009   : cube_lut_0 = 14'b10100000011110;
        10'd1010   : cube_lut_0 = 14'b10100000100010;
        10'd1011   : cube_lut_0 = 14'b10100000100101;
        10'd1012   : cube_lut_0 = 14'b10100000101000;
        10'd1013   : cube_lut_0 = 14'b10100000101100;
        10'd1014   : cube_lut_0 = 14'b10100000101111;
        10'd1015   : cube_lut_0 = 14'b10100000110010;
        10'd1016   : cube_lut_0 = 14'b10100000110110;
        10'd1017   : cube_lut_0 = 14'b10100000111001;
        10'd1018   : cube_lut_0 = 14'b10100000111101;
        10'd1019   : cube_lut_0 = 14'b10100001000000;
        10'd1020   : cube_lut_0 = 14'b10100001000011;
        10'd1021   : cube_lut_0 = 14'b10100001000111;
        10'd1022   : cube_lut_0 = 14'b10100001001010;
        10'd1023   : cube_lut_0 = 14'b10100001001101;
        
        
    endcase
end

always@* begin
    
    cube_lut_1 = 0;
    
    case(i_data[9:0])
        
        10'd0   : cube_lut_1    = 14'b10100001010001;
        10'd1   : cube_lut_1    = 14'b10100001010100;
        10'd2   : cube_lut_1    = 14'b10100001010111;
        10'd3   : cube_lut_1    = 14'b10100001011011;
        10'd4   : cube_lut_1    = 14'b10100001011110;
        10'd5   : cube_lut_1    = 14'b10100001100010;
        10'd6   : cube_lut_1    = 14'b10100001100101;
        10'd7   : cube_lut_1    = 14'b10100001101000;
        10'd8   : cube_lut_1    = 14'b10100001101100;
        10'd9   : cube_lut_1    = 14'b10100001101111;
        10'd10   : cube_lut_1   = 14'b10100001110010;
        10'd11   : cube_lut_1   = 14'b10100001110110;
        10'd12   : cube_lut_1   = 14'b10100001111001;
        10'd13   : cube_lut_1   = 14'b10100001111100;
        10'd14   : cube_lut_1   = 14'b10100010000000;
        10'd15   : cube_lut_1   = 14'b10100010000011;
        10'd16   : cube_lut_1   = 14'b10100010000110;
        10'd17   : cube_lut_1   = 14'b10100010001010;
        10'd18   : cube_lut_1   = 14'b10100010001101;
        10'd19   : cube_lut_1   = 14'b10100010010000;
        10'd20   : cube_lut_1   = 14'b10100010010100;
        10'd21   : cube_lut_1   = 14'b10100010010111;
        10'd22   : cube_lut_1   = 14'b10100010011010;
        10'd23   : cube_lut_1   = 14'b10100010011101;
        10'd24   : cube_lut_1   = 14'b10100010100001;
        10'd25   : cube_lut_1   = 14'b10100010100100;
        10'd26   : cube_lut_1   = 14'b10100010100111;
        10'd27   : cube_lut_1   = 14'b10100010101011;
        10'd28   : cube_lut_1   = 14'b10100010101110;
        10'd29   : cube_lut_1   = 14'b10100010110001;
        10'd30   : cube_lut_1   = 14'b10100010110101;
        10'd31   : cube_lut_1   = 14'b10100010111000;
        10'd32   : cube_lut_1   = 14'b10100010111011;
        10'd33   : cube_lut_1   = 14'b10100010111110;
        10'd34   : cube_lut_1   = 14'b10100011000010;
        10'd35   : cube_lut_1   = 14'b10100011000101;
        10'd36   : cube_lut_1   = 14'b10100011001000;
        10'd37   : cube_lut_1   = 14'b10100011001100;
        10'd38   : cube_lut_1   = 14'b10100011001111;
        10'd39   : cube_lut_1   = 14'b10100011010010;
        10'd40   : cube_lut_1   = 14'b10100011010101;
        10'd41   : cube_lut_1   = 14'b10100011011001;
        10'd42   : cube_lut_1   = 14'b10100011011100;
        10'd43   : cube_lut_1   = 14'b10100011011111;
        10'd44   : cube_lut_1   = 14'b10100011100011;
        10'd45   : cube_lut_1   = 14'b10100011100110;
        10'd46   : cube_lut_1   = 14'b10100011101001;
        10'd47   : cube_lut_1   = 14'b10100011101100;
        10'd48   : cube_lut_1   = 14'b10100011110000;
        10'd49   : cube_lut_1   = 14'b10100011110011;
        10'd50   : cube_lut_1   = 14'b10100011110110;
        10'd51   : cube_lut_1   = 14'b10100011111001;
        10'd52   : cube_lut_1   = 14'b10100011111101;
        10'd53   : cube_lut_1   = 14'b10100100000000;
        10'd54   : cube_lut_1   = 14'b10100100000011;
        10'd55   : cube_lut_1   = 14'b10100100000110;
        10'd56   : cube_lut_1   = 14'b10100100001010;
        10'd57   : cube_lut_1   = 14'b10100100001101;
        10'd58   : cube_lut_1   = 14'b10100100010000;
        10'd59   : cube_lut_1   = 14'b10100100010011;
        10'd60   : cube_lut_1   = 14'b10100100010111;
        10'd61   : cube_lut_1   = 14'b10100100011010;
        10'd62   : cube_lut_1   = 14'b10100100011101;
        10'd63   : cube_lut_1   = 14'b10100100100000;
        10'd64   : cube_lut_1   = 14'b10100100100011;
        10'd65   : cube_lut_1   = 14'b10100100100111;
        10'd66   : cube_lut_1   = 14'b10100100101010;
        10'd67   : cube_lut_1   = 14'b10100100101101;
        10'd68   : cube_lut_1   = 14'b10100100110000;
        10'd69   : cube_lut_1   = 14'b10100100110100;
        10'd70   : cube_lut_1   = 14'b10100100110111;
        10'd71   : cube_lut_1   = 14'b10100100111010;
        10'd72   : cube_lut_1   = 14'b10100100111101;
        10'd73   : cube_lut_1   = 14'b10100101000000;
        10'd74   : cube_lut_1   = 14'b10100101000100;
        10'd75   : cube_lut_1   = 14'b10100101000111;
        10'd76   : cube_lut_1   = 14'b10100101001010;
        10'd77   : cube_lut_1   = 14'b10100101001101;
        10'd78   : cube_lut_1   = 14'b10100101010000;
        10'd79   : cube_lut_1   = 14'b10100101010100;
        10'd80   : cube_lut_1   = 14'b10100101010111;
        10'd81   : cube_lut_1   = 14'b10100101011010;
        10'd82   : cube_lut_1   = 14'b10100101011101;
        10'd83   : cube_lut_1   = 14'b10100101100000;
        10'd84   : cube_lut_1   = 14'b10100101100100;
        10'd85   : cube_lut_1   = 14'b10100101100111;
        10'd86   : cube_lut_1   = 14'b10100101101010;
        10'd87   : cube_lut_1   = 14'b10100101101101;
        10'd88   : cube_lut_1   = 14'b10100101110000;
        10'd89   : cube_lut_1   = 14'b10100101110100;
        10'd90   : cube_lut_1   = 14'b10100101110111;
        10'd91   : cube_lut_1   = 14'b10100101111010;
        10'd92   : cube_lut_1   = 14'b10100101111101;
        10'd93   : cube_lut_1   = 14'b10100110000000;
        10'd94   : cube_lut_1   = 14'b10100110000011;
        10'd95   : cube_lut_1   = 14'b10100110000111;
        10'd96   : cube_lut_1   = 14'b10100110001010;
        10'd97   : cube_lut_1   = 14'b10100110001101;
        10'd98   : cube_lut_1   = 14'b10100110010000;
        10'd99   : cube_lut_1   = 14'b10100110010011;
        10'd100   : cube_lut_1  = 14'b10100110010110;
        10'd101   : cube_lut_1  = 14'b10100110011010;
        10'd102   : cube_lut_1  = 14'b10100110011101;
        10'd103   : cube_lut_1  = 14'b10100110100000;
        10'd104   : cube_lut_1  = 14'b10100110100011;
        10'd105   : cube_lut_1  = 14'b10100110100110;
        10'd106   : cube_lut_1  = 14'b10100110101001;
        10'd107   : cube_lut_1  = 14'b10100110101100;
        10'd108   : cube_lut_1  = 14'b10100110110000;
        10'd109   : cube_lut_1  = 14'b10100110110011;
        10'd110   : cube_lut_1  = 14'b10100110110110;
        10'd111   : cube_lut_1  = 14'b10100110111001;
        10'd112   : cube_lut_1  = 14'b10100110111100;
        10'd113   : cube_lut_1  = 14'b10100110111111;
        10'd114   : cube_lut_1  = 14'b10100111000010;
        10'd115   : cube_lut_1  = 14'b10100111000110;
        10'd116   : cube_lut_1  = 14'b10100111001001;
        10'd117   : cube_lut_1  = 14'b10100111001100;
        10'd118   : cube_lut_1  = 14'b10100111001111;
        10'd119   : cube_lut_1  = 14'b10100111010010;
        10'd120   : cube_lut_1  = 14'b10100111010101;
        10'd121   : cube_lut_1  = 14'b10100111011000;
        10'd122   : cube_lut_1  = 14'b10100111011011;
        10'd123   : cube_lut_1  = 14'b10100111011111;
        10'd124   : cube_lut_1  = 14'b10100111100010;
        10'd125   : cube_lut_1  = 14'b10100111100101;
        10'd126   : cube_lut_1  = 14'b10100111101000;
        10'd127   : cube_lut_1  = 14'b10100111101011;
        10'd128   : cube_lut_1  = 14'b10100111101110;
        10'd129   : cube_lut_1  = 14'b10100111110001;
        10'd130   : cube_lut_1  = 14'b10100111110100;
        10'd131   : cube_lut_1  = 14'b10100111110111;
        10'd132   : cube_lut_1  = 14'b10100111111010;
        10'd133   : cube_lut_1  = 14'b10100111111110;
        10'd134   : cube_lut_1  = 14'b10101000000001;
        10'd135   : cube_lut_1  = 14'b10101000000100;
        10'd136   : cube_lut_1  = 14'b10101000000111;
        10'd137   : cube_lut_1  = 14'b10101000001010;
        10'd138   : cube_lut_1  = 14'b10101000001101;
        10'd139   : cube_lut_1  = 14'b10101000010000;
        10'd140   : cube_lut_1  = 14'b10101000010011;
        10'd141   : cube_lut_1  = 14'b10101000010110;
        10'd142   : cube_lut_1  = 14'b10101000011001;
        10'd143   : cube_lut_1  = 14'b10101000011100;
        10'd144   : cube_lut_1  = 14'b10101000100000;
        10'd145   : cube_lut_1  = 14'b10101000100011;
        10'd146   : cube_lut_1  = 14'b10101000100110;
        10'd147   : cube_lut_1  = 14'b10101000101001;
        10'd148   : cube_lut_1  = 14'b10101000101100;
        10'd149   : cube_lut_1  = 14'b10101000101111;
        10'd150   : cube_lut_1  = 14'b10101000110010;
        10'd151   : cube_lut_1  = 14'b10101000110101;
        10'd152   : cube_lut_1  = 14'b10101000111000;
        10'd153   : cube_lut_1  = 14'b10101000111011;
        10'd154   : cube_lut_1  = 14'b10101000111110;
        10'd155   : cube_lut_1  = 14'b10101001000001;
        10'd156   : cube_lut_1  = 14'b10101001000100;
        10'd157   : cube_lut_1  = 14'b10101001000111;
        10'd158   : cube_lut_1  = 14'b10101001001010;
        10'd159   : cube_lut_1  = 14'b10101001001101;
        10'd160   : cube_lut_1  = 14'b10101001010001;
        10'd161   : cube_lut_1  = 14'b10101001010100;
        10'd162   : cube_lut_1  = 14'b10101001010111;
        10'd163   : cube_lut_1  = 14'b10101001011010;
        10'd164   : cube_lut_1  = 14'b10101001011101;
        10'd165   : cube_lut_1  = 14'b10101001100000;
        10'd166   : cube_lut_1  = 14'b10101001100011;
        10'd167   : cube_lut_1  = 14'b10101001100110;
        10'd168   : cube_lut_1  = 14'b10101001101001;
        10'd169   : cube_lut_1  = 14'b10101001101100;
        10'd170   : cube_lut_1  = 14'b10101001101111;
        10'd171   : cube_lut_1  = 14'b10101001110010;
        10'd172   : cube_lut_1  = 14'b10101001110101;
        10'd173   : cube_lut_1  = 14'b10101001111000;
        10'd174   : cube_lut_1  = 14'b10101001111011;
        10'd175   : cube_lut_1  = 14'b10101001111110;
        10'd176   : cube_lut_1  = 14'b10101010000001;
        10'd177   : cube_lut_1  = 14'b10101010000100;
        10'd178   : cube_lut_1  = 14'b10101010000111;
        10'd179   : cube_lut_1  = 14'b10101010001010;
        10'd180   : cube_lut_1  = 14'b10101010001101;
        10'd181   : cube_lut_1  = 14'b10101010010000;
        10'd182   : cube_lut_1  = 14'b10101010010011;
        10'd183   : cube_lut_1  = 14'b10101010010110;
        10'd184   : cube_lut_1  = 14'b10101010011001;
        10'd185   : cube_lut_1  = 14'b10101010011100;
        10'd186   : cube_lut_1  = 14'b10101010011111;
        10'd187   : cube_lut_1  = 14'b10101010100010;
        10'd188   : cube_lut_1  = 14'b10101010100101;
        10'd189   : cube_lut_1  = 14'b10101010101000;
        10'd190   : cube_lut_1  = 14'b10101010101011;
        10'd191   : cube_lut_1  = 14'b10101010101110;
        10'd192   : cube_lut_1  = 14'b10101010110001;
        10'd193   : cube_lut_1  = 14'b10101010110100;
        10'd194   : cube_lut_1  = 14'b10101010110111;
        10'd195   : cube_lut_1  = 14'b10101010111010;
        10'd196   : cube_lut_1  = 14'b10101010111101;
        10'd197   : cube_lut_1  = 14'b10101011000000;
        10'd198   : cube_lut_1  = 14'b10101011000011;
        10'd199   : cube_lut_1  = 14'b10101011000110;
        10'd200   : cube_lut_1  = 14'b10101011001001;
        10'd201   : cube_lut_1  = 14'b10101011001100;
        10'd202   : cube_lut_1  = 14'b10101011001111;
        10'd203   : cube_lut_1  = 14'b10101011010010;
        10'd204   : cube_lut_1  = 14'b10101011010101;
        10'd205   : cube_lut_1  = 14'b10101011011000;
        10'd206   : cube_lut_1  = 14'b10101011011011;
        10'd207   : cube_lut_1  = 14'b10101011011110;
        10'd208   : cube_lut_1  = 14'b10101011100001;
        10'd209   : cube_lut_1  = 14'b10101011100100;
        10'd210   : cube_lut_1  = 14'b10101011100111;
        10'd211   : cube_lut_1  = 14'b10101011101010;
        10'd212   : cube_lut_1  = 14'b10101011101101;
        10'd213   : cube_lut_1  = 14'b10101011110000;
        10'd214   : cube_lut_1  = 14'b10101011110011;
        10'd215   : cube_lut_1  = 14'b10101011110110;
        10'd216   : cube_lut_1  = 14'b10101011111001;
        10'd217   : cube_lut_1  = 14'b10101011111100;
        10'd218   : cube_lut_1  = 14'b10101011111111;
        10'd219   : cube_lut_1  = 14'b10101100000010;
        10'd220   : cube_lut_1  = 14'b10101100000101;
        10'd221   : cube_lut_1  = 14'b10101100000111;
        10'd222   : cube_lut_1  = 14'b10101100001010;
        10'd223   : cube_lut_1  = 14'b10101100001101;
        10'd224   : cube_lut_1  = 14'b10101100010000;
        10'd225   : cube_lut_1  = 14'b10101100010011;
        10'd226   : cube_lut_1  = 14'b10101100010110;
        10'd227   : cube_lut_1  = 14'b10101100011001;
        10'd228   : cube_lut_1  = 14'b10101100011100;
        10'd229   : cube_lut_1  = 14'b10101100011111;
        10'd230   : cube_lut_1  = 14'b10101100100010;
        10'd231   : cube_lut_1  = 14'b10101100100101;
        10'd232   : cube_lut_1  = 14'b10101100101000;
        10'd233   : cube_lut_1  = 14'b10101100101011;
        10'd234   : cube_lut_1  = 14'b10101100101110;
        10'd235   : cube_lut_1  = 14'b10101100110001;
        10'd236   : cube_lut_1  = 14'b10101100110100;
        10'd237   : cube_lut_1  = 14'b10101100110110;
        10'd238   : cube_lut_1  = 14'b10101100111001;
        10'd239   : cube_lut_1  = 14'b10101100111100;
        10'd240   : cube_lut_1  = 14'b10101100111111;
        10'd241   : cube_lut_1  = 14'b10101101000010;
        10'd242   : cube_lut_1  = 14'b10101101000101;
        10'd243   : cube_lut_1  = 14'b10101101001000;
        10'd244   : cube_lut_1  = 14'b10101101001011;
        10'd245   : cube_lut_1  = 14'b10101101001110;
        10'd246   : cube_lut_1  = 14'b10101101010001;
        10'd247   : cube_lut_1  = 14'b10101101010100;
        10'd248   : cube_lut_1  = 14'b10101101010111;
        10'd249   : cube_lut_1  = 14'b10101101011001;
        10'd250   : cube_lut_1  = 14'b10101101011100;
        10'd251   : cube_lut_1  = 14'b10101101011111;
        10'd252   : cube_lut_1  = 14'b10101101100010;
        10'd253   : cube_lut_1  = 14'b10101101100101;
        10'd254   : cube_lut_1  = 14'b10101101101000;
        10'd255   : cube_lut_1  = 14'b10101101101011;
        10'd256   : cube_lut_1  = 14'b10101101101110;
        10'd257   : cube_lut_1  = 14'b10101101110001;
        10'd258   : cube_lut_1  = 14'b10101101110100;
        10'd259   : cube_lut_1  = 14'b10101101110110;
        10'd260   : cube_lut_1  = 14'b10101101111001;
        10'd261   : cube_lut_1  = 14'b10101101111100;
        10'd262   : cube_lut_1  = 14'b10101101111111;
        10'd263   : cube_lut_1  = 14'b10101110000010;
        10'd264   : cube_lut_1  = 14'b10101110000101;
        10'd265   : cube_lut_1  = 14'b10101110001000;
        10'd266   : cube_lut_1  = 14'b10101110001011;
        10'd267   : cube_lut_1  = 14'b10101110001110;
        10'd268   : cube_lut_1  = 14'b10101110010000;
        10'd269   : cube_lut_1  = 14'b10101110010011;
        10'd270   : cube_lut_1  = 14'b10101110010110;
        10'd271   : cube_lut_1  = 14'b10101110011001;
        10'd272   : cube_lut_1  = 14'b10101110011100;
        10'd273   : cube_lut_1  = 14'b10101110011111;
        10'd274   : cube_lut_1  = 14'b10101110100010;
        10'd275   : cube_lut_1  = 14'b10101110100100;
        10'd276   : cube_lut_1  = 14'b10101110100111;
        10'd277   : cube_lut_1  = 14'b10101110101010;
        10'd278   : cube_lut_1  = 14'b10101110101101;
        10'd279   : cube_lut_1  = 14'b10101110110000;
        10'd280   : cube_lut_1  = 14'b10101110110011;
        10'd281   : cube_lut_1  = 14'b10101110110110;
        10'd282   : cube_lut_1  = 14'b10101110111001;
        10'd283   : cube_lut_1  = 14'b10101110111011;
        10'd284   : cube_lut_1  = 14'b10101110111110;
        10'd285   : cube_lut_1  = 14'b10101111000001;
        10'd286   : cube_lut_1  = 14'b10101111000100;
        10'd287   : cube_lut_1  = 14'b10101111000111;
        10'd288   : cube_lut_1  = 14'b10101111001010;
        10'd289   : cube_lut_1  = 14'b10101111001100;
        10'd290   : cube_lut_1  = 14'b10101111001111;
        10'd291   : cube_lut_1  = 14'b10101111010010;
        10'd292   : cube_lut_1  = 14'b10101111010101;
        10'd293   : cube_lut_1  = 14'b10101111011000;
        10'd294   : cube_lut_1  = 14'b10101111011011;
        10'd295   : cube_lut_1  = 14'b10101111011110;
        10'd296   : cube_lut_1  = 14'b10101111100000;
        10'd297   : cube_lut_1  = 14'b10101111100011;
        10'd298   : cube_lut_1  = 14'b10101111100110;
        10'd299   : cube_lut_1  = 14'b10101111101001;
        10'd300   : cube_lut_1  = 14'b10101111101100;
        10'd301   : cube_lut_1  = 14'b10101111101111;
        10'd302   : cube_lut_1  = 14'b10101111110001;
        10'd303   : cube_lut_1  = 14'b10101111110100;
        10'd304   : cube_lut_1  = 14'b10101111110111;
        10'd305   : cube_lut_1  = 14'b10101111111010;
        10'd306   : cube_lut_1  = 14'b10101111111101;
        10'd307   : cube_lut_1  = 14'b10110000000000;
        10'd308   : cube_lut_1  = 14'b10110000000010;
        10'd309   : cube_lut_1  = 14'b10110000000101;
        10'd310   : cube_lut_1  = 14'b10110000001000;
        10'd311   : cube_lut_1  = 14'b10110000001011;
        10'd312   : cube_lut_1  = 14'b10110000001110;
        10'd313   : cube_lut_1  = 14'b10110000010000;
        10'd314   : cube_lut_1  = 14'b10110000010011;
        10'd315   : cube_lut_1  = 14'b10110000010110;
        10'd316   : cube_lut_1  = 14'b10110000011001;
        10'd317   : cube_lut_1  = 14'b10110000011100;
        10'd318   : cube_lut_1  = 14'b10110000011110;
        10'd319   : cube_lut_1  = 14'b10110000100001;
        10'd320   : cube_lut_1  = 14'b10110000100100;
        10'd321   : cube_lut_1  = 14'b10110000100111;
        10'd322   : cube_lut_1  = 14'b10110000101010;
        10'd323   : cube_lut_1  = 14'b10110000101100;
        10'd324   : cube_lut_1  = 14'b10110000101111;
        10'd325   : cube_lut_1  = 14'b10110000110010;
        10'd326   : cube_lut_1  = 14'b10110000110101;
        10'd327   : cube_lut_1  = 14'b10110000111000;
        10'd328   : cube_lut_1  = 14'b10110000111010;
        10'd329   : cube_lut_1  = 14'b10110000111101;
        10'd330   : cube_lut_1  = 14'b10110001000000;
        10'd331   : cube_lut_1  = 14'b10110001000011;
        10'd332   : cube_lut_1  = 14'b10110001000110;
        10'd333   : cube_lut_1  = 14'b10110001001000;
        10'd334   : cube_lut_1  = 14'b10110001001011;
        10'd335   : cube_lut_1  = 14'b10110001001110;
        10'd336   : cube_lut_1  = 14'b10110001010001;
        10'd337   : cube_lut_1  = 14'b10110001010100;
        10'd338   : cube_lut_1  = 14'b10110001010110;
        10'd339   : cube_lut_1  = 14'b10110001011001;
        10'd340   : cube_lut_1  = 14'b10110001011100;
        10'd341   : cube_lut_1  = 14'b10110001011111;
        10'd342   : cube_lut_1  = 14'b10110001100001;
        10'd343   : cube_lut_1  = 14'b10110001100100;
        10'd344   : cube_lut_1  = 14'b10110001100111;
        10'd345   : cube_lut_1  = 14'b10110001101010;
        10'd346   : cube_lut_1  = 14'b10110001101100;
        10'd347   : cube_lut_1  = 14'b10110001101111;
        10'd348   : cube_lut_1  = 14'b10110001110010;
        10'd349   : cube_lut_1  = 14'b10110001110101;
        10'd350   : cube_lut_1  = 14'b10110001111000;
        10'd351   : cube_lut_1  = 14'b10110001111010;
        10'd352   : cube_lut_1  = 14'b10110001111101;
        10'd353   : cube_lut_1  = 14'b10110010000000;
        10'd354   : cube_lut_1  = 14'b10110010000011;
        10'd355   : cube_lut_1  = 14'b10110010000101;
        10'd356   : cube_lut_1  = 14'b10110010001000;
        10'd357   : cube_lut_1  = 14'b10110010001011;
        10'd358   : cube_lut_1  = 14'b10110010001110;
        10'd359   : cube_lut_1  = 14'b10110010010000;
        10'd360   : cube_lut_1  = 14'b10110010010011;
        10'd361   : cube_lut_1  = 14'b10110010010110;
        10'd362   : cube_lut_1  = 14'b10110010011001;
        10'd363   : cube_lut_1  = 14'b10110010011011;
        10'd364   : cube_lut_1  = 14'b10110010011110;
        10'd365   : cube_lut_1  = 14'b10110010100001;
        10'd366   : cube_lut_1  = 14'b10110010100100;
        10'd367   : cube_lut_1  = 14'b10110010100110;
        10'd368   : cube_lut_1  = 14'b10110010101001;
        10'd369   : cube_lut_1  = 14'b10110010101100;
        10'd370   : cube_lut_1  = 14'b10110010101110;
        10'd371   : cube_lut_1  = 14'b10110010110001;
        10'd372   : cube_lut_1  = 14'b10110010110100;
        10'd373   : cube_lut_1  = 14'b10110010110111;
        10'd374   : cube_lut_1  = 14'b10110010111001;
        10'd375   : cube_lut_1  = 14'b10110010111100;
        10'd376   : cube_lut_1  = 14'b10110010111111;
        10'd377   : cube_lut_1  = 14'b10110011000010;
        10'd378   : cube_lut_1  = 14'b10110011000100;
        10'd379   : cube_lut_1  = 14'b10110011000111;
        10'd380   : cube_lut_1  = 14'b10110011001010;
        10'd381   : cube_lut_1  = 14'b10110011001100;
        10'd382   : cube_lut_1  = 14'b10110011001111;
        10'd383   : cube_lut_1  = 14'b10110011010010;
        10'd384   : cube_lut_1  = 14'b10110011010101;
        10'd385   : cube_lut_1  = 14'b10110011010111;
        10'd386   : cube_lut_1  = 14'b10110011011010;
        10'd387   : cube_lut_1  = 14'b10110011011101;
        10'd388   : cube_lut_1  = 14'b10110011100000;
        10'd389   : cube_lut_1  = 14'b10110011100010;
        10'd390   : cube_lut_1  = 14'b10110011100101;
        10'd391   : cube_lut_1  = 14'b10110011101000;
        10'd392   : cube_lut_1  = 14'b10110011101010;
        10'd393   : cube_lut_1  = 14'b10110011101101;
        10'd394   : cube_lut_1  = 14'b10110011110000;
        10'd395   : cube_lut_1  = 14'b10110011110010;
        10'd396   : cube_lut_1  = 14'b10110011110101;
        10'd397   : cube_lut_1  = 14'b10110011111000;
        10'd398   : cube_lut_1  = 14'b10110011111011;
        10'd399   : cube_lut_1  = 14'b10110011111101;
        10'd400   : cube_lut_1  = 14'b10110100000000;
        10'd401   : cube_lut_1  = 14'b10110100000011;
        10'd402   : cube_lut_1  = 14'b10110100000101;
        10'd403   : cube_lut_1  = 14'b10110100001000;
        10'd404   : cube_lut_1  = 14'b10110100001011;
        10'd405   : cube_lut_1  = 14'b10110100001101;
        10'd406   : cube_lut_1  = 14'b10110100010000;
        10'd407   : cube_lut_1  = 14'b10110100010011;
        10'd408   : cube_lut_1  = 14'b10110100010101;
        10'd409   : cube_lut_1  = 14'b10110100011000;
        10'd410   : cube_lut_1  = 14'b10110100011011;
        10'd411   : cube_lut_1  = 14'b10110100011110;
        10'd412   : cube_lut_1  = 14'b10110100100000;
        10'd413   : cube_lut_1  = 14'b10110100100011;
        10'd414   : cube_lut_1  = 14'b10110100100110;
        10'd415   : cube_lut_1  = 14'b10110100101000;
        10'd416   : cube_lut_1  = 14'b10110100101011;
        10'd417   : cube_lut_1  = 14'b10110100101110;
        10'd418   : cube_lut_1  = 14'b10110100110000;
        10'd419   : cube_lut_1  = 14'b10110100110011;
        10'd420   : cube_lut_1  = 14'b10110100110110;
        10'd421   : cube_lut_1  = 14'b10110100111000;
        10'd422   : cube_lut_1  = 14'b10110100111011;
        10'd423   : cube_lut_1  = 14'b10110100111110;
        10'd424   : cube_lut_1  = 14'b10110101000000;
        10'd425   : cube_lut_1  = 14'b10110101000011;
        10'd426   : cube_lut_1  = 14'b10110101000110;
        10'd427   : cube_lut_1  = 14'b10110101001000;
        10'd428   : cube_lut_1  = 14'b10110101001011;
        10'd429   : cube_lut_1  = 14'b10110101001110;
        10'd430   : cube_lut_1  = 14'b10110101010000;
        10'd431   : cube_lut_1  = 14'b10110101010011;
        10'd432   : cube_lut_1  = 14'b10110101010110;
        10'd433   : cube_lut_1  = 14'b10110101011000;
        10'd434   : cube_lut_1  = 14'b10110101011011;
        10'd435   : cube_lut_1  = 14'b10110101011110;
        10'd436   : cube_lut_1  = 14'b10110101100000;
        10'd437   : cube_lut_1  = 14'b10110101100011;
        10'd438   : cube_lut_1  = 14'b10110101100110;
        10'd439   : cube_lut_1  = 14'b10110101101000;
        10'd440   : cube_lut_1  = 14'b10110101101011;
        10'd441   : cube_lut_1  = 14'b10110101101101;
        10'd442   : cube_lut_1  = 14'b10110101110000;
        10'd443   : cube_lut_1  = 14'b10110101110011;
        10'd444   : cube_lut_1  = 14'b10110101110101;
        10'd445   : cube_lut_1  = 14'b10110101111000;
        10'd446   : cube_lut_1  = 14'b10110101111011;
        10'd447   : cube_lut_1  = 14'b10110101111101;
        10'd448   : cube_lut_1  = 14'b10110110000000;
        10'd449   : cube_lut_1  = 14'b10110110000011;
        10'd450   : cube_lut_1  = 14'b10110110000101;
        10'd451   : cube_lut_1  = 14'b10110110001000;
        10'd452   : cube_lut_1  = 14'b10110110001011;
        10'd453   : cube_lut_1  = 14'b10110110001101;
        10'd454   : cube_lut_1  = 14'b10110110010000;
        10'd455   : cube_lut_1  = 14'b10110110010010;
        10'd456   : cube_lut_1  = 14'b10110110010101;
        10'd457   : cube_lut_1  = 14'b10110110011000;
        10'd458   : cube_lut_1  = 14'b10110110011010;
        10'd459   : cube_lut_1  = 14'b10110110011101;
        10'd460   : cube_lut_1  = 14'b10110110100000;
        10'd461   : cube_lut_1  = 14'b10110110100010;
        10'd462   : cube_lut_1  = 14'b10110110100101;
        10'd463   : cube_lut_1  = 14'b10110110100111;
        10'd464   : cube_lut_1  = 14'b10110110101010;
        10'd465   : cube_lut_1  = 14'b10110110101101;
        10'd466   : cube_lut_1  = 14'b10110110101111;
        10'd467   : cube_lut_1  = 14'b10110110110010;
        10'd468   : cube_lut_1  = 14'b10110110110100;
        10'd469   : cube_lut_1  = 14'b10110110110111;
        10'd470   : cube_lut_1  = 14'b10110110111010;
        10'd471   : cube_lut_1  = 14'b10110110111100;
        10'd472   : cube_lut_1  = 14'b10110110111111;
        10'd473   : cube_lut_1  = 14'b10110111000010;
        10'd474   : cube_lut_1  = 14'b10110111000100;
        10'd475   : cube_lut_1  = 14'b10110111000111;
        10'd476   : cube_lut_1  = 14'b10110111001001;
        10'd477   : cube_lut_1  = 14'b10110111001100;
        10'd478   : cube_lut_1  = 14'b10110111001111;
        10'd479   : cube_lut_1  = 14'b10110111010001;
        10'd480   : cube_lut_1  = 14'b10110111010100;
        10'd481   : cube_lut_1  = 14'b10110111010110;
        10'd482   : cube_lut_1  = 14'b10110111011001;
        10'd483   : cube_lut_1  = 14'b10110111011100;
        10'd484   : cube_lut_1  = 14'b10110111011110;
        10'd485   : cube_lut_1  = 14'b10110111100001;
        10'd486   : cube_lut_1  = 14'b10110111100011;
        10'd487   : cube_lut_1  = 14'b10110111100110;
        10'd488   : cube_lut_1  = 14'b10110111101001;
        10'd489   : cube_lut_1  = 14'b10110111101011;
        10'd490   : cube_lut_1  = 14'b10110111101110;
        10'd491   : cube_lut_1  = 14'b10110111110000;
        10'd492   : cube_lut_1  = 14'b10110111110011;
        10'd493   : cube_lut_1  = 14'b10110111110101;
        10'd494   : cube_lut_1  = 14'b10110111111000;
        10'd495   : cube_lut_1  = 14'b10110111111011;
        10'd496   : cube_lut_1  = 14'b10110111111101;
        10'd497   : cube_lut_1  = 14'b10111000000000;
        10'd498   : cube_lut_1  = 14'b10111000000010;
        10'd499   : cube_lut_1  = 14'b10111000000101;
        10'd500   : cube_lut_1  = 14'b10111000001000;
        10'd501   : cube_lut_1  = 14'b10111000001010;
        10'd502   : cube_lut_1  = 14'b10111000001101;
        10'd503   : cube_lut_1  = 14'b10111000001111;
        10'd504   : cube_lut_1  = 14'b10111000010010;
        10'd505   : cube_lut_1  = 14'b10111000010100;
        10'd506   : cube_lut_1  = 14'b10111000010111;
        10'd507   : cube_lut_1  = 14'b10111000011010;
        10'd508   : cube_lut_1  = 14'b10111000011100;
        10'd509   : cube_lut_1  = 14'b10111000011111;
        10'd510   : cube_lut_1  = 14'b10111000100001;
        10'd511   : cube_lut_1  = 14'b10111000100100;
        10'd512   : cube_lut_1  = 14'b10111000100110;
        10'd513   : cube_lut_1  = 14'b10111000101001;
        10'd514   : cube_lut_1  = 14'b10111000101100;
        10'd515   : cube_lut_1  = 14'b10111000101110;
        10'd516   : cube_lut_1  = 14'b10111000110001;
        10'd517   : cube_lut_1  = 14'b10111000110011;
        10'd518   : cube_lut_1  = 14'b10111000110110;
        10'd519   : cube_lut_1  = 14'b10111000111000;
        10'd520   : cube_lut_1  = 14'b10111000111011;
        10'd521   : cube_lut_1  = 14'b10111000111101;
        10'd522   : cube_lut_1  = 14'b10111001000000;
        10'd523   : cube_lut_1  = 14'b10111001000011;
        10'd524   : cube_lut_1  = 14'b10111001000101;
        10'd525   : cube_lut_1  = 14'b10111001001000;
        10'd526   : cube_lut_1  = 14'b10111001001010;
        10'd527   : cube_lut_1  = 14'b10111001001101;
        10'd528   : cube_lut_1  = 14'b10111001001111;
        10'd529   : cube_lut_1  = 14'b10111001010010;
        10'd530   : cube_lut_1  = 14'b10111001010100;
        10'd531   : cube_lut_1  = 14'b10111001010111;
        10'd532   : cube_lut_1  = 14'b10111001011001;
        10'd533   : cube_lut_1  = 14'b10111001011100;
        10'd534   : cube_lut_1  = 14'b10111001011111;
        10'd535   : cube_lut_1  = 14'b10111001100001;
        10'd536   : cube_lut_1  = 14'b10111001100100;
        10'd537   : cube_lut_1  = 14'b10111001100110;
        10'd538   : cube_lut_1  = 14'b10111001101001;
        10'd539   : cube_lut_1  = 14'b10111001101011;
        10'd540   : cube_lut_1  = 14'b10111001101110;
        10'd541   : cube_lut_1  = 14'b10111001110000;
        10'd542   : cube_lut_1  = 14'b10111001110011;
        10'd543   : cube_lut_1  = 14'b10111001110101;
        10'd544   : cube_lut_1  = 14'b10111001111000;
        10'd545   : cube_lut_1  = 14'b10111001111010;
        10'd546   : cube_lut_1  = 14'b10111001111101;
        10'd547   : cube_lut_1  = 14'b10111001111111;
        10'd548   : cube_lut_1  = 14'b10111010000010;
        10'd549   : cube_lut_1  = 14'b10111010000101;
        10'd550   : cube_lut_1  = 14'b10111010000111;
        10'd551   : cube_lut_1  = 14'b10111010001010;
        10'd552   : cube_lut_1  = 14'b10111010001100;
        10'd553   : cube_lut_1  = 14'b10111010001111;
        10'd554   : cube_lut_1  = 14'b10111010010001;
        10'd555   : cube_lut_1  = 14'b10111010010100;
        10'd556   : cube_lut_1  = 14'b10111010010110;
        10'd557   : cube_lut_1  = 14'b10111010011001;
        10'd558   : cube_lut_1  = 14'b10111010011011;
        10'd559   : cube_lut_1  = 14'b10111010011110;
        10'd560   : cube_lut_1  = 14'b10111010100000;
        10'd561   : cube_lut_1  = 14'b10111010100011;
        10'd562   : cube_lut_1  = 14'b10111010100101;
        10'd563   : cube_lut_1  = 14'b10111010101000;
        10'd564   : cube_lut_1  = 14'b10111010101010;
        10'd565   : cube_lut_1  = 14'b10111010101101;
        10'd566   : cube_lut_1  = 14'b10111010101111;
        10'd567   : cube_lut_1  = 14'b10111010110010;
        10'd568   : cube_lut_1  = 14'b10111010110100;
        10'd569   : cube_lut_1  = 14'b10111010110111;
        10'd570   : cube_lut_1  = 14'b10111010111001;
        10'd571   : cube_lut_1  = 14'b10111010111100;
        10'd572   : cube_lut_1  = 14'b10111010111110;
        10'd573   : cube_lut_1  = 14'b10111011000001;
        10'd574   : cube_lut_1  = 14'b10111011000011;
        10'd575   : cube_lut_1  = 14'b10111011000110;
        10'd576   : cube_lut_1  = 14'b10111011001000;
        10'd577   : cube_lut_1  = 14'b10111011001011;
        10'd578   : cube_lut_1  = 14'b10111011001101;
        10'd579   : cube_lut_1  = 14'b10111011010000;
        10'd580   : cube_lut_1  = 14'b10111011010010;
        10'd581   : cube_lut_1  = 14'b10111011010101;
        10'd582   : cube_lut_1  = 14'b10111011010111;
        10'd583   : cube_lut_1  = 14'b10111011011010;
        10'd584   : cube_lut_1  = 14'b10111011011100;
        10'd585   : cube_lut_1  = 14'b10111011011111;
        10'd586   : cube_lut_1  = 14'b10111011100001;
        10'd587   : cube_lut_1  = 14'b10111011100100;
        10'd588   : cube_lut_1  = 14'b10111011100110;
        10'd589   : cube_lut_1  = 14'b10111011101001;
        10'd590   : cube_lut_1  = 14'b10111011101011;
        10'd591   : cube_lut_1  = 14'b10111011101110;
        10'd592   : cube_lut_1  = 14'b10111011110000;
        10'd593   : cube_lut_1  = 14'b10111011110011;
        10'd594   : cube_lut_1  = 14'b10111011110101;
        10'd595   : cube_lut_1  = 14'b10111011110111;
        10'd596   : cube_lut_1  = 14'b10111011111010;
        10'd597   : cube_lut_1  = 14'b10111011111100;
        10'd598   : cube_lut_1  = 14'b10111011111111;
        10'd599   : cube_lut_1  = 14'b10111100000001;
        10'd600   : cube_lut_1  = 14'b10111100000100;
        10'd601   : cube_lut_1  = 14'b10111100000110;
        10'd602   : cube_lut_1  = 14'b10111100001001;
        10'd603   : cube_lut_1  = 14'b10111100001011;
        10'd604   : cube_lut_1  = 14'b10111100001110;
        10'd605   : cube_lut_1  = 14'b10111100010000;
        10'd606   : cube_lut_1  = 14'b10111100010011;
        10'd607   : cube_lut_1  = 14'b10111100010101;
        10'd608   : cube_lut_1  = 14'b10111100011000;
        10'd609   : cube_lut_1  = 14'b10111100011010;
        10'd610   : cube_lut_1  = 14'b10111100011101;
        10'd611   : cube_lut_1  = 14'b10111100011111;
        10'd612   : cube_lut_1  = 14'b10111100100001;
        10'd613   : cube_lut_1  = 14'b10111100100100;
        10'd614   : cube_lut_1  = 14'b10111100100110;
        10'd615   : cube_lut_1  = 14'b10111100101001;
        10'd616   : cube_lut_1  = 14'b10111100101011;
        10'd617   : cube_lut_1  = 14'b10111100101110;
        10'd618   : cube_lut_1  = 14'b10111100110000;
        10'd619   : cube_lut_1  = 14'b10111100110011;
        10'd620   : cube_lut_1  = 14'b10111100110101;
        10'd621   : cube_lut_1  = 14'b10111100111000;
        10'd622   : cube_lut_1  = 14'b10111100111010;
        10'd623   : cube_lut_1  = 14'b10111100111100;
        10'd624   : cube_lut_1  = 14'b10111100111111;
        10'd625   : cube_lut_1  = 14'b10111101000001;
        10'd626   : cube_lut_1  = 14'b10111101000100;
        10'd627   : cube_lut_1  = 14'b10111101000110;
        10'd628   : cube_lut_1  = 14'b10111101001001;
        10'd629   : cube_lut_1  = 14'b10111101001011;
        10'd630   : cube_lut_1  = 14'b10111101001110;
        10'd631   : cube_lut_1  = 14'b10111101010000;
        10'd632   : cube_lut_1  = 14'b10111101010010;
        10'd633   : cube_lut_1  = 14'b10111101010101;
        10'd634   : cube_lut_1  = 14'b10111101010111;
        10'd635   : cube_lut_1  = 14'b10111101011010;
        10'd636   : cube_lut_1  = 14'b10111101011100;
        10'd637   : cube_lut_1  = 14'b10111101011111;
        10'd638   : cube_lut_1  = 14'b10111101100001;
        10'd639   : cube_lut_1  = 14'b10111101100011;
        10'd640   : cube_lut_1  = 14'b10111101100110;
        10'd641   : cube_lut_1  = 14'b10111101101000;
        10'd642   : cube_lut_1  = 14'b10111101101011;
        10'd643   : cube_lut_1  = 14'b10111101101101;
        10'd644   : cube_lut_1  = 14'b10111101110000;
        10'd645   : cube_lut_1  = 14'b10111101110010;
        10'd646   : cube_lut_1  = 14'b10111101110100;
        10'd647   : cube_lut_1  = 14'b10111101110111;
        10'd648   : cube_lut_1  = 14'b10111101111001;
        10'd649   : cube_lut_1  = 14'b10111101111100;
        10'd650   : cube_lut_1  = 14'b10111101111110;
        10'd651   : cube_lut_1  = 14'b10111110000001;
        10'd652   : cube_lut_1  = 14'b10111110000011;
        10'd653   : cube_lut_1  = 14'b10111110000101;
        10'd654   : cube_lut_1  = 14'b10111110001000;
        10'd655   : cube_lut_1  = 14'b10111110001010;
        10'd656   : cube_lut_1  = 14'b10111110001101;
        10'd657   : cube_lut_1  = 14'b10111110001111;
        10'd658   : cube_lut_1  = 14'b10111110010001;
        10'd659   : cube_lut_1  = 14'b10111110010100;
        10'd660   : cube_lut_1  = 14'b10111110010110;
        10'd661   : cube_lut_1  = 14'b10111110011001;
        10'd662   : cube_lut_1  = 14'b10111110011011;
        10'd663   : cube_lut_1  = 14'b10111110011110;
        10'd664   : cube_lut_1  = 14'b10111110100000;
        10'd665   : cube_lut_1  = 14'b10111110100010;
        10'd666   : cube_lut_1  = 14'b10111110100101;
        10'd667   : cube_lut_1  = 14'b10111110100111;
        10'd668   : cube_lut_1  = 14'b10111110101010;
        10'd669   : cube_lut_1  = 14'b10111110101100;
        10'd670   : cube_lut_1  = 14'b10111110101110;
        10'd671   : cube_lut_1  = 14'b10111110110001;
        10'd672   : cube_lut_1  = 14'b10111110110011;
        10'd673   : cube_lut_1  = 14'b10111110110110;
        10'd674   : cube_lut_1  = 14'b10111110111000;
        10'd675   : cube_lut_1  = 14'b10111110111010;
        10'd676   : cube_lut_1  = 14'b10111110111101;
        10'd677   : cube_lut_1  = 14'b10111110111111;
        10'd678   : cube_lut_1  = 14'b10111111000010;
        10'd679   : cube_lut_1  = 14'b10111111000100;
        10'd680   : cube_lut_1  = 14'b10111111000110;
        10'd681   : cube_lut_1  = 14'b10111111001001;
        10'd682   : cube_lut_1  = 14'b10111111001011;
        10'd683   : cube_lut_1  = 14'b10111111001110;
        10'd684   : cube_lut_1  = 14'b10111111010000;
        10'd685   : cube_lut_1  = 14'b10111111010010;
        10'd686   : cube_lut_1  = 14'b10111111010101;
        10'd687   : cube_lut_1  = 14'b10111111010111;
        10'd688   : cube_lut_1  = 14'b10111111011001;
        10'd689   : cube_lut_1  = 14'b10111111011100;
        10'd690   : cube_lut_1  = 14'b10111111011110;
        10'd691   : cube_lut_1  = 14'b10111111100001;
        10'd692   : cube_lut_1  = 14'b10111111100011;
        10'd693   : cube_lut_1  = 14'b10111111100101;
        10'd694   : cube_lut_1  = 14'b10111111101000;
        10'd695   : cube_lut_1  = 14'b10111111101010;
        10'd696   : cube_lut_1  = 14'b10111111101101;
        10'd697   : cube_lut_1  = 14'b10111111101111;
        10'd698   : cube_lut_1  = 14'b10111111110001;
        10'd699   : cube_lut_1  = 14'b10111111110100;
        10'd700   : cube_lut_1  = 14'b10111111110110;
        10'd701   : cube_lut_1  = 14'b10111111111000;
        10'd702   : cube_lut_1  = 14'b10111111111011;
        10'd703   : cube_lut_1  = 14'b10111111111101;
        10'd704   : cube_lut_1  = 14'b11000000000000;
        10'd705   : cube_lut_1  = 14'b11000000000010;
        10'd706   : cube_lut_1  = 14'b11000000000100;
        10'd707   : cube_lut_1  = 14'b11000000000111;
        10'd708   : cube_lut_1  = 14'b11000000001001;
        10'd709   : cube_lut_1  = 14'b11000000001011;
        10'd710   : cube_lut_1  = 14'b11000000001110;
        10'd711   : cube_lut_1  = 14'b11000000010000;
        10'd712   : cube_lut_1  = 14'b11000000010010;
        10'd713   : cube_lut_1  = 14'b11000000010101;
        10'd714   : cube_lut_1  = 14'b11000000010111;
        10'd715   : cube_lut_1  = 14'b11000000011010;
        10'd716   : cube_lut_1  = 14'b11000000011100;
        10'd717   : cube_lut_1  = 14'b11000000011110;
        10'd718   : cube_lut_1  = 14'b11000000100001;
        10'd719   : cube_lut_1  = 14'b11000000100011;
        10'd720   : cube_lut_1  = 14'b11000000100101;
        10'd721   : cube_lut_1  = 14'b11000000101000;
        10'd722   : cube_lut_1  = 14'b11000000101010;
        10'd723   : cube_lut_1  = 14'b11000000101100;
        10'd724   : cube_lut_1  = 14'b11000000101111;
        10'd725   : cube_lut_1  = 14'b11000000110001;
        10'd726   : cube_lut_1  = 14'b11000000110011;
        10'd727   : cube_lut_1  = 14'b11000000110110;
        10'd728   : cube_lut_1  = 14'b11000000111000;
        10'd729   : cube_lut_1  = 14'b11000000111010;
        10'd730   : cube_lut_1  = 14'b11000000111101;
        10'd731   : cube_lut_1  = 14'b11000000111111;
        10'd732   : cube_lut_1  = 14'b11000001000010;
        10'd733   : cube_lut_1  = 14'b11000001000100;
        10'd734   : cube_lut_1  = 14'b11000001000110;
        10'd735   : cube_lut_1  = 14'b11000001001001;
        10'd736   : cube_lut_1  = 14'b11000001001011;
        10'd737   : cube_lut_1  = 14'b11000001001101;
        10'd738   : cube_lut_1  = 14'b11000001010000;
        10'd739   : cube_lut_1  = 14'b11000001010010;
        10'd740   : cube_lut_1  = 14'b11000001010100;
        10'd741   : cube_lut_1  = 14'b11000001010111;
        10'd742   : cube_lut_1  = 14'b11000001011001;
        10'd743   : cube_lut_1  = 14'b11000001011011;
        10'd744   : cube_lut_1  = 14'b11000001011110;
        10'd745   : cube_lut_1  = 14'b11000001100000;
        10'd746   : cube_lut_1  = 14'b11000001100010;
        10'd747   : cube_lut_1  = 14'b11000001100101;
        10'd748   : cube_lut_1  = 14'b11000001100111;
        10'd749   : cube_lut_1  = 14'b11000001101001;
        10'd750   : cube_lut_1  = 14'b11000001101100;
        10'd751   : cube_lut_1  = 14'b11000001101110;
        10'd752   : cube_lut_1  = 14'b11000001110000;
        10'd753   : cube_lut_1  = 14'b11000001110011;
        10'd754   : cube_lut_1  = 14'b11000001110101;
        10'd755   : cube_lut_1  = 14'b11000001110111;
        10'd756   : cube_lut_1  = 14'b11000001111010;
        10'd757   : cube_lut_1  = 14'b11000001111100;
        10'd758   : cube_lut_1  = 14'b11000001111110;
        10'd759   : cube_lut_1  = 14'b11000010000001;
        10'd760   : cube_lut_1  = 14'b11000010000011;
        10'd761   : cube_lut_1  = 14'b11000010000101;
        10'd762   : cube_lut_1  = 14'b11000010000111;
        10'd763   : cube_lut_1  = 14'b11000010001010;
        10'd764   : cube_lut_1  = 14'b11000010001100;
        10'd765   : cube_lut_1  = 14'b11000010001110;
        10'd766   : cube_lut_1  = 14'b11000010010001;
        10'd767   : cube_lut_1  = 14'b11000010010011;
        10'd768   : cube_lut_1  = 14'b11000010010101;
        10'd769   : cube_lut_1  = 14'b11000010011000;
        10'd770   : cube_lut_1  = 14'b11000010011010;
        10'd771   : cube_lut_1  = 14'b11000010011100;
        10'd772   : cube_lut_1  = 14'b11000010011111;
        10'd773   : cube_lut_1  = 14'b11000010100001;
        10'd774   : cube_lut_1  = 14'b11000010100011;
        10'd775   : cube_lut_1  = 14'b11000010100110;
        10'd776   : cube_lut_1  = 14'b11000010101000;
        10'd777   : cube_lut_1  = 14'b11000010101010;
        10'd778   : cube_lut_1  = 14'b11000010101100;
        10'd779   : cube_lut_1  = 14'b11000010101111;
        10'd780   : cube_lut_1  = 14'b11000010110001;
        10'd781   : cube_lut_1  = 14'b11000010110011;
        10'd782   : cube_lut_1  = 14'b11000010110110;
        10'd783   : cube_lut_1  = 14'b11000010111000;
        10'd784   : cube_lut_1  = 14'b11000010111010;
        10'd785   : cube_lut_1  = 14'b11000010111101;
        10'd786   : cube_lut_1  = 14'b11000010111111;
        10'd787   : cube_lut_1  = 14'b11000011000001;
        10'd788   : cube_lut_1  = 14'b11000011000011;
        10'd789   : cube_lut_1  = 14'b11000011000110;
        10'd790   : cube_lut_1  = 14'b11000011001000;
        10'd791   : cube_lut_1  = 14'b11000011001010;
        10'd792   : cube_lut_1  = 14'b11000011001101;
        10'd793   : cube_lut_1  = 14'b11000011001111;
        10'd794   : cube_lut_1  = 14'b11000011010001;
        10'd795   : cube_lut_1  = 14'b11000011010100;
        10'd796   : cube_lut_1  = 14'b11000011010110;
        10'd797   : cube_lut_1  = 14'b11000011011000;
        10'd798   : cube_lut_1  = 14'b11000011011010;
        10'd799   : cube_lut_1  = 14'b11000011011101;
        10'd800   : cube_lut_1  = 14'b11000011011111;
        10'd801   : cube_lut_1  = 14'b11000011100001;
        10'd802   : cube_lut_1  = 14'b11000011100100;
        10'd803   : cube_lut_1  = 14'b11000011100110;
        10'd804   : cube_lut_1  = 14'b11000011101000;
        10'd805   : cube_lut_1  = 14'b11000011101010;
        10'd806   : cube_lut_1  = 14'b11000011101101;
        10'd807   : cube_lut_1  = 14'b11000011101111;
        10'd808   : cube_lut_1  = 14'b11000011110001;
        10'd809   : cube_lut_1  = 14'b11000011110100;
        10'd810   : cube_lut_1  = 14'b11000011110110;
        10'd811   : cube_lut_1  = 14'b11000011111000;
        10'd812   : cube_lut_1  = 14'b11000011111010;
        10'd813   : cube_lut_1  = 14'b11000011111101;
        10'd814   : cube_lut_1  = 14'b11000011111111;
        10'd815   : cube_lut_1  = 14'b11000100000001;
        10'd816   : cube_lut_1  = 14'b11000100000011;
        10'd817   : cube_lut_1  = 14'b11000100000110;
        10'd818   : cube_lut_1  = 14'b11000100001000;
        10'd819   : cube_lut_1  = 14'b11000100001010;
        10'd820   : cube_lut_1  = 14'b11000100001101;
        10'd821   : cube_lut_1  = 14'b11000100001111;
        10'd822   : cube_lut_1  = 14'b11000100010001;
        10'd823   : cube_lut_1  = 14'b11000100010011;
        10'd824   : cube_lut_1  = 14'b11000100010110;
        10'd825   : cube_lut_1  = 14'b11000100011000;
        10'd826   : cube_lut_1  = 14'b11000100011010;
        10'd827   : cube_lut_1  = 14'b11000100011100;
        10'd828   : cube_lut_1  = 14'b11000100011111;
        10'd829   : cube_lut_1  = 14'b11000100100001;
        10'd830   : cube_lut_1  = 14'b11000100100011;
        10'd831   : cube_lut_1  = 14'b11000100100101;
        10'd832   : cube_lut_1  = 14'b11000100101000;
        10'd833   : cube_lut_1  = 14'b11000100101010;
        10'd834   : cube_lut_1  = 14'b11000100101100;
        10'd835   : cube_lut_1  = 14'b11000100101110;
        10'd836   : cube_lut_1  = 14'b11000100110001;
        10'd837   : cube_lut_1  = 14'b11000100110011;
        10'd838   : cube_lut_1  = 14'b11000100110101;
        10'd839   : cube_lut_1  = 14'b11000100111000;
        10'd840   : cube_lut_1  = 14'b11000100111010;
        10'd841   : cube_lut_1  = 14'b11000100111100;
        10'd842   : cube_lut_1  = 14'b11000100111110;
        10'd843   : cube_lut_1  = 14'b11000101000001;
        10'd844   : cube_lut_1  = 14'b11000101000011;
        10'd845   : cube_lut_1  = 14'b11000101000101;
        10'd846   : cube_lut_1  = 14'b11000101000111;
        10'd847   : cube_lut_1  = 14'b11000101001010;
        10'd848   : cube_lut_1  = 14'b11000101001100;
        10'd849   : cube_lut_1  = 14'b11000101001110;
        10'd850   : cube_lut_1  = 14'b11000101010000;
        10'd851   : cube_lut_1  = 14'b11000101010011;
        10'd852   : cube_lut_1  = 14'b11000101010101;
        10'd853   : cube_lut_1  = 14'b11000101010111;
        10'd854   : cube_lut_1  = 14'b11000101011001;
        10'd855   : cube_lut_1  = 14'b11000101011011;
        10'd856   : cube_lut_1  = 14'b11000101011110;
        10'd857   : cube_lut_1  = 14'b11000101100000;
        10'd858   : cube_lut_1  = 14'b11000101100010;
        10'd859   : cube_lut_1  = 14'b11000101100100;
        10'd860   : cube_lut_1  = 14'b11000101100111;
        10'd861   : cube_lut_1  = 14'b11000101101001;
        10'd862   : cube_lut_1  = 14'b11000101101011;
        10'd863   : cube_lut_1  = 14'b11000101101101;
        10'd864   : cube_lut_1  = 14'b11000101110000;
        10'd865   : cube_lut_1  = 14'b11000101110010;
        10'd866   : cube_lut_1  = 14'b11000101110100;
        10'd867   : cube_lut_1  = 14'b11000101110110;
        10'd868   : cube_lut_1  = 14'b11000101111001;
        10'd869   : cube_lut_1  = 14'b11000101111011;
        10'd870   : cube_lut_1  = 14'b11000101111101;
        10'd871   : cube_lut_1  = 14'b11000101111111;
        10'd872   : cube_lut_1  = 14'b11000110000001;
        10'd873   : cube_lut_1  = 14'b11000110000100;
        10'd874   : cube_lut_1  = 14'b11000110000110;
        10'd875   : cube_lut_1  = 14'b11000110001000;
        10'd876   : cube_lut_1  = 14'b11000110001010;
        10'd877   : cube_lut_1  = 14'b11000110001101;
        10'd878   : cube_lut_1  = 14'b11000110001111;
        10'd879   : cube_lut_1  = 14'b11000110010001;
        10'd880   : cube_lut_1  = 14'b11000110010011;
        10'd881   : cube_lut_1  = 14'b11000110010101;
        10'd882   : cube_lut_1  = 14'b11000110011000;
        10'd883   : cube_lut_1  = 14'b11000110011010;
        10'd884   : cube_lut_1  = 14'b11000110011100;
        10'd885   : cube_lut_1  = 14'b11000110011110;
        10'd886   : cube_lut_1  = 14'b11000110100001;
        10'd887   : cube_lut_1  = 14'b11000110100011;
        10'd888   : cube_lut_1  = 14'b11000110100101;
        10'd889   : cube_lut_1  = 14'b11000110100111;
        10'd890   : cube_lut_1  = 14'b11000110101001;
        10'd891   : cube_lut_1  = 14'b11000110101100;
        10'd892   : cube_lut_1  = 14'b11000110101110;
        10'd893   : cube_lut_1  = 14'b11000110110000;
        10'd894   : cube_lut_1  = 14'b11000110110010;
        10'd895   : cube_lut_1  = 14'b11000110110101;
        10'd896   : cube_lut_1  = 14'b11000110110111;
        10'd897   : cube_lut_1  = 14'b11000110111001;
        10'd898   : cube_lut_1  = 14'b11000110111011;
        10'd899   : cube_lut_1  = 14'b11000110111101;
        10'd900   : cube_lut_1  = 14'b11000111000000;
        10'd901   : cube_lut_1  = 14'b11000111000010;
        10'd902   : cube_lut_1  = 14'b11000111000100;
        10'd903   : cube_lut_1  = 14'b11000111000110;
        10'd904   : cube_lut_1  = 14'b11000111001000;
        10'd905   : cube_lut_1  = 14'b11000111001011;
        10'd906   : cube_lut_1  = 14'b11000111001101;
        10'd907   : cube_lut_1  = 14'b11000111001111;
        10'd908   : cube_lut_1  = 14'b11000111010001;
        10'd909   : cube_lut_1  = 14'b11000111010011;
        10'd910   : cube_lut_1  = 14'b11000111010110;
        10'd911   : cube_lut_1  = 14'b11000111011000;
        10'd912   : cube_lut_1  = 14'b11000111011010;
        10'd913   : cube_lut_1  = 14'b11000111011100;
        10'd914   : cube_lut_1  = 14'b11000111011110;
        10'd915   : cube_lut_1  = 14'b11000111100001;
        10'd916   : cube_lut_1  = 14'b11000111100011;
        10'd917   : cube_lut_1  = 14'b11000111100101;
        10'd918   : cube_lut_1  = 14'b11000111100111;
        10'd919   : cube_lut_1  = 14'b11000111101001;
        10'd920   : cube_lut_1  = 14'b11000111101100;
        10'd921   : cube_lut_1  = 14'b11000111101110;
        10'd922   : cube_lut_1  = 14'b11000111110000;
        10'd923   : cube_lut_1  = 14'b11000111110010;
        10'd924   : cube_lut_1  = 14'b11000111110100;
        10'd925   : cube_lut_1  = 14'b11000111110110;
        10'd926   : cube_lut_1  = 14'b11000111111001;
        10'd927   : cube_lut_1  = 14'b11000111111011;
        10'd928   : cube_lut_1  = 14'b11000111111101;
        10'd929   : cube_lut_1  = 14'b11000111111111;
        10'd930   : cube_lut_1  = 14'b11001000000001;
        10'd931   : cube_lut_1  = 14'b11001000000100;
        10'd932   : cube_lut_1  = 14'b11001000000110;
        10'd933   : cube_lut_1  = 14'b11001000001000;
        10'd934   : cube_lut_1  = 14'b11001000001010;
        10'd935   : cube_lut_1  = 14'b11001000001100;
        10'd936   : cube_lut_1  = 14'b11001000001111;
        10'd937   : cube_lut_1  = 14'b11001000010001;
        10'd938   : cube_lut_1  = 14'b11001000010011;
        10'd939   : cube_lut_1  = 14'b11001000010101;
        10'd940   : cube_lut_1  = 14'b11001000010111;
        10'd941   : cube_lut_1  = 14'b11001000011001;
        10'd942   : cube_lut_1  = 14'b11001000011100;
        10'd943   : cube_lut_1  = 14'b11001000011110;
        10'd944   : cube_lut_1  = 14'b11001000100000;
        10'd945   : cube_lut_1  = 14'b11001000100010;
        10'd946   : cube_lut_1  = 14'b11001000100100;
        10'd947   : cube_lut_1  = 14'b11001000100110;
        10'd948   : cube_lut_1  = 14'b11001000101001;
        10'd949   : cube_lut_1  = 14'b11001000101011;
        10'd950   : cube_lut_1  = 14'b11001000101101;
        10'd951   : cube_lut_1  = 14'b11001000101111;
        10'd952   : cube_lut_1  = 14'b11001000110001;
        10'd953   : cube_lut_1  = 14'b11001000110011;
        10'd954   : cube_lut_1  = 14'b11001000110110;
        10'd955   : cube_lut_1  = 14'b11001000111000;
        10'd956   : cube_lut_1  = 14'b11001000111010;
        10'd957   : cube_lut_1  = 14'b11001000111100;
        10'd958   : cube_lut_1  = 14'b11001000111110;
        10'd959   : cube_lut_1  = 14'b11001001000000;
        10'd960   : cube_lut_1  = 14'b11001001000011;
        10'd961   : cube_lut_1  = 14'b11001001000101;
        10'd962   : cube_lut_1  = 14'b11001001000111;
        10'd963   : cube_lut_1  = 14'b11001001001001;
        10'd964   : cube_lut_1  = 14'b11001001001011;
        10'd965   : cube_lut_1  = 14'b11001001001101;
        10'd966   : cube_lut_1  = 14'b11001001010000;
        10'd967   : cube_lut_1  = 14'b11001001010010;
        10'd968   : cube_lut_1  = 14'b11001001010100;
        10'd969   : cube_lut_1  = 14'b11001001010110;
        10'd970   : cube_lut_1  = 14'b11001001011000;
        10'd971   : cube_lut_1  = 14'b11001001011010;
        10'd972   : cube_lut_1  = 14'b11001001011100;
        10'd973   : cube_lut_1  = 14'b11001001011111;
        10'd974   : cube_lut_1  = 14'b11001001100001;
        10'd975   : cube_lut_1  = 14'b11001001100011;
        10'd976   : cube_lut_1  = 14'b11001001100101;
        10'd977   : cube_lut_1  = 14'b11001001100111;
        10'd978   : cube_lut_1  = 14'b11001001101001;
        10'd979   : cube_lut_1  = 14'b11001001101100;
        10'd980   : cube_lut_1  = 14'b11001001101110;
        10'd981   : cube_lut_1  = 14'b11001001110000;
        10'd982   : cube_lut_1  = 14'b11001001110010;
        10'd983   : cube_lut_1  = 14'b11001001110100;
        10'd984   : cube_lut_1  = 14'b11001001110110;
        10'd985   : cube_lut_1  = 14'b11001001111000;
        10'd986   : cube_lut_1  = 14'b11001001111011;
        10'd987   : cube_lut_1  = 14'b11001001111101;
        10'd988   : cube_lut_1  = 14'b11001001111111;
        10'd989   : cube_lut_1  = 14'b11001010000001;
        10'd990   : cube_lut_1  = 14'b11001010000011;
        10'd991   : cube_lut_1  = 14'b11001010000101;
        10'd992   : cube_lut_1  = 14'b11001010000111;
        10'd993   : cube_lut_1  = 14'b11001010001010;
        10'd994   : cube_lut_1  = 14'b11001010001100;
        10'd995   : cube_lut_1  = 14'b11001010001110;
        10'd996   : cube_lut_1  = 14'b11001010010000;
        10'd997   : cube_lut_1  = 14'b11001010010010;
        10'd998   : cube_lut_1  = 14'b11001010010100;
        10'd999   : cube_lut_1  = 14'b11001010010110;
        10'd1000   : cube_lut_1 = 14'b11001010011000;
        10'd1001   : cube_lut_1 = 14'b11001010011011;
        10'd1002   : cube_lut_1 = 14'b11001010011101;
        10'd1003   : cube_lut_1 = 14'b11001010011111;
        10'd1004   : cube_lut_1 = 14'b11001010100001;
        10'd1005   : cube_lut_1 = 14'b11001010100011;
        10'd1006   : cube_lut_1 = 14'b11001010100101;
        10'd1007   : cube_lut_1 = 14'b11001010100111;
        10'd1008   : cube_lut_1 = 14'b11001010101010;
        10'd1009   : cube_lut_1 = 14'b11001010101100;
        10'd1010   : cube_lut_1 = 14'b11001010101110;
        10'd1011   : cube_lut_1 = 14'b11001010110000;
        10'd1012   : cube_lut_1 = 14'b11001010110010;
        10'd1013   : cube_lut_1 = 14'b11001010110100;
        10'd1014   : cube_lut_1 = 14'b11001010110110;
        10'd1015   : cube_lut_1 = 14'b11001010111000;
        10'd1016   : cube_lut_1 = 14'b11001010111011;
        10'd1017   : cube_lut_1 = 14'b11001010111101;
        10'd1018   : cube_lut_1 = 14'b11001010111111;
        10'd1019   : cube_lut_1 = 14'b11001011000001;
        10'd1020   : cube_lut_1 = 14'b11001011000011;
        10'd1021   : cube_lut_1 = 14'b11001011000101;
        10'd1022   : cube_lut_1 = 14'b11001011000111;
        10'd1023   : cube_lut_1 = 14'b11001011001001;
        
    endcase
end

always@* begin
    
    cube_lut_2 = 0;
    
    case(i_data[9:0])
        
        10'd0   : cube_lut_2    = 14'b11001011001011;
        10'd1   : cube_lut_2    = 14'b11001011001110;
        10'd2   : cube_lut_2    = 14'b11001011010000;
        10'd3   : cube_lut_2    = 14'b11001011010010;
        10'd4   : cube_lut_2    = 14'b11001011010100;
        10'd5   : cube_lut_2    = 14'b11001011010110;
        10'd6   : cube_lut_2    = 14'b11001011011000;
        10'd7   : cube_lut_2    = 14'b11001011011010;
        10'd8   : cube_lut_2    = 14'b11001011011100;
        10'd9   : cube_lut_2    = 14'b11001011011111;
        10'd10   : cube_lut_2   = 14'b11001011100001;
        10'd11   : cube_lut_2   = 14'b11001011100011;
        10'd12   : cube_lut_2   = 14'b11001011100101;
        10'd13   : cube_lut_2   = 14'b11001011100111;
        10'd14   : cube_lut_2   = 14'b11001011101001;
        10'd15   : cube_lut_2   = 14'b11001011101011;
        10'd16   : cube_lut_2   = 14'b11001011101101;
        10'd17   : cube_lut_2   = 14'b11001011101111;
        10'd18   : cube_lut_2   = 14'b11001011110001;
        10'd19   : cube_lut_2   = 14'b11001011110100;
        10'd20   : cube_lut_2   = 14'b11001011110110;
        10'd21   : cube_lut_2   = 14'b11001011111000;
        10'd22   : cube_lut_2   = 14'b11001011111010;
        10'd23   : cube_lut_2   = 14'b11001011111100;
        10'd24   : cube_lut_2   = 14'b11001011111110;
        10'd25   : cube_lut_2   = 14'b11001100000000;
        10'd26   : cube_lut_2   = 14'b11001100000010;
        10'd27   : cube_lut_2   = 14'b11001100000100;
        10'd28   : cube_lut_2   = 14'b11001100000110;
        10'd29   : cube_lut_2   = 14'b11001100001001;
        10'd30   : cube_lut_2   = 14'b11001100001011;
        10'd31   : cube_lut_2   = 14'b11001100001101;
        10'd32   : cube_lut_2   = 14'b11001100001111;
        10'd33   : cube_lut_2   = 14'b11001100010001;
        10'd34   : cube_lut_2   = 14'b11001100010011;
        10'd35   : cube_lut_2   = 14'b11001100010101;
        10'd36   : cube_lut_2   = 14'b11001100010111;
        10'd37   : cube_lut_2   = 14'b11001100011001;
        10'd38   : cube_lut_2   = 14'b11001100011011;
        10'd39   : cube_lut_2   = 14'b11001100011110;
        10'd40   : cube_lut_2   = 14'b11001100100000;
        10'd41   : cube_lut_2   = 14'b11001100100010;
        10'd42   : cube_lut_2   = 14'b11001100100100;
        10'd43   : cube_lut_2   = 14'b11001100100110;
        10'd44   : cube_lut_2   = 14'b11001100101000;
        10'd45   : cube_lut_2   = 14'b11001100101010;
        10'd46   : cube_lut_2   = 14'b11001100101100;
        10'd47   : cube_lut_2   = 14'b11001100101110;
        10'd48   : cube_lut_2   = 14'b11001100110000;
        10'd49   : cube_lut_2   = 14'b11001100110010;
        10'd50   : cube_lut_2   = 14'b11001100110100;
        10'd51   : cube_lut_2   = 14'b11001100110111;
        10'd52   : cube_lut_2   = 14'b11001100111001;
        10'd53   : cube_lut_2   = 14'b11001100111011;
        10'd54   : cube_lut_2   = 14'b11001100111101;
        10'd55   : cube_lut_2   = 14'b11001100111111;
        10'd56   : cube_lut_2   = 14'b11001101000001;
        10'd57   : cube_lut_2   = 14'b11001101000011;
        10'd58   : cube_lut_2   = 14'b11001101000101;
        10'd59   : cube_lut_2   = 14'b11001101000111;
        10'd60   : cube_lut_2   = 14'b11001101001001;
        10'd61   : cube_lut_2   = 14'b11001101001011;
        10'd62   : cube_lut_2   = 14'b11001101001101;
        10'd63   : cube_lut_2   = 14'b11001101001111;
        10'd64   : cube_lut_2   = 14'b11001101010010;
        10'd65   : cube_lut_2   = 14'b11001101010100;
        10'd66   : cube_lut_2   = 14'b11001101010110;
        10'd67   : cube_lut_2   = 14'b11001101011000;
        10'd68   : cube_lut_2   = 14'b11001101011010;
        10'd69   : cube_lut_2   = 14'b11001101011100;
        10'd70   : cube_lut_2   = 14'b11001101011110;
        10'd71   : cube_lut_2   = 14'b11001101100000;
        10'd72   : cube_lut_2   = 14'b11001101100010;
        10'd73   : cube_lut_2   = 14'b11001101100100;
        10'd74   : cube_lut_2   = 14'b11001101100110;
        10'd75   : cube_lut_2   = 14'b11001101101000;
        10'd76   : cube_lut_2   = 14'b11001101101010;
        10'd77   : cube_lut_2   = 14'b11001101101100;
        10'd78   : cube_lut_2   = 14'b11001101101111;
        10'd79   : cube_lut_2   = 14'b11001101110001;
        10'd80   : cube_lut_2   = 14'b11001101110011;
        10'd81   : cube_lut_2   = 14'b11001101110101;
        10'd82   : cube_lut_2   = 14'b11001101110111;
        10'd83   : cube_lut_2   = 14'b11001101111001;
        10'd84   : cube_lut_2   = 14'b11001101111011;
        10'd85   : cube_lut_2   = 14'b11001101111101;
        10'd86   : cube_lut_2   = 14'b11001101111111;
        10'd87   : cube_lut_2   = 14'b11001110000001;
        10'd88   : cube_lut_2   = 14'b11001110000011;
        10'd89   : cube_lut_2   = 14'b11001110000101;
        10'd90   : cube_lut_2   = 14'b11001110000111;
        10'd91   : cube_lut_2   = 14'b11001110001001;
        10'd92   : cube_lut_2   = 14'b11001110001011;
        10'd93   : cube_lut_2   = 14'b11001110001101;
        10'd94   : cube_lut_2   = 14'b11001110001111;
        10'd95   : cube_lut_2   = 14'b11001110010010;
        10'd96   : cube_lut_2   = 14'b11001110010100;
        10'd97   : cube_lut_2   = 14'b11001110010110;
        10'd98   : cube_lut_2   = 14'b11001110011000;
        10'd99   : cube_lut_2   = 14'b11001110011010;
        10'd100   : cube_lut_2  = 14'b11001110011100;
        10'd101   : cube_lut_2  = 14'b11001110011110;
        10'd102   : cube_lut_2  = 14'b11001110100000;
        10'd103   : cube_lut_2  = 14'b11001110100010;
        10'd104   : cube_lut_2  = 14'b11001110100100;
        10'd105   : cube_lut_2  = 14'b11001110100110;
        10'd106   : cube_lut_2  = 14'b11001110101000;
        10'd107   : cube_lut_2  = 14'b11001110101010;
        10'd108   : cube_lut_2  = 14'b11001110101100;
        10'd109   : cube_lut_2  = 14'b11001110101110;
        10'd110   : cube_lut_2  = 14'b11001110110000;
        10'd111   : cube_lut_2  = 14'b11001110110010;
        10'd112   : cube_lut_2  = 14'b11001110110100;
        10'd113   : cube_lut_2  = 14'b11001110110110;
        10'd114   : cube_lut_2  = 14'b11001110111000;
        10'd115   : cube_lut_2  = 14'b11001110111010;
        10'd116   : cube_lut_2  = 14'b11001110111101;
        10'd117   : cube_lut_2  = 14'b11001110111111;
        10'd118   : cube_lut_2  = 14'b11001111000001;
        10'd119   : cube_lut_2  = 14'b11001111000011;
        10'd120   : cube_lut_2  = 14'b11001111000101;
        10'd121   : cube_lut_2  = 14'b11001111000111;
        10'd122   : cube_lut_2  = 14'b11001111001001;
        10'd123   : cube_lut_2  = 14'b11001111001011;
        10'd124   : cube_lut_2  = 14'b11001111001101;
        10'd125   : cube_lut_2  = 14'b11001111001111;
        10'd126   : cube_lut_2  = 14'b11001111010001;
        10'd127   : cube_lut_2  = 14'b11001111010011;
        10'd128   : cube_lut_2  = 14'b11001111010101;
        10'd129   : cube_lut_2  = 14'b11001111010111;
        10'd130   : cube_lut_2  = 14'b11001111011001;
        10'd131   : cube_lut_2  = 14'b11001111011011;
        10'd132   : cube_lut_2  = 14'b11001111011101;
        10'd133   : cube_lut_2  = 14'b11001111011111;
        10'd134   : cube_lut_2  = 14'b11001111100001;
        10'd135   : cube_lut_2  = 14'b11001111100011;
        10'd136   : cube_lut_2  = 14'b11001111100101;
        10'd137   : cube_lut_2  = 14'b11001111100111;
        10'd138   : cube_lut_2  = 14'b11001111101001;
        10'd139   : cube_lut_2  = 14'b11001111101011;
        10'd140   : cube_lut_2  = 14'b11001111101101;
        10'd141   : cube_lut_2  = 14'b11001111101111;
        10'd142   : cube_lut_2  = 14'b11001111110001;
        10'd143   : cube_lut_2  = 14'b11001111110011;
        10'd144   : cube_lut_2  = 14'b11001111110101;
        10'd145   : cube_lut_2  = 14'b11001111110111;
        10'd146   : cube_lut_2  = 14'b11001111111001;
        10'd147   : cube_lut_2  = 14'b11001111111011;
        10'd148   : cube_lut_2  = 14'b11001111111101;
        10'd149   : cube_lut_2  = 14'b11010000000000;
        10'd150   : cube_lut_2  = 14'b11010000000010;
        10'd151   : cube_lut_2  = 14'b11010000000100;
        10'd152   : cube_lut_2  = 14'b11010000000110;
        10'd153   : cube_lut_2  = 14'b11010000001000;
        10'd154   : cube_lut_2  = 14'b11010000001010;
        10'd155   : cube_lut_2  = 14'b11010000001100;
        10'd156   : cube_lut_2  = 14'b11010000001110;
        10'd157   : cube_lut_2  = 14'b11010000010000;
        10'd158   : cube_lut_2  = 14'b11010000010010;
        10'd159   : cube_lut_2  = 14'b11010000010100;
        10'd160   : cube_lut_2  = 14'b11010000010110;
        10'd161   : cube_lut_2  = 14'b11010000011000;
        10'd162   : cube_lut_2  = 14'b11010000011010;
        10'd163   : cube_lut_2  = 14'b11010000011100;
        10'd164   : cube_lut_2  = 14'b11010000011110;
        10'd165   : cube_lut_2  = 14'b11010000100000;
        10'd166   : cube_lut_2  = 14'b11010000100010;
        10'd167   : cube_lut_2  = 14'b11010000100100;
        10'd168   : cube_lut_2  = 14'b11010000100110;
        10'd169   : cube_lut_2  = 14'b11010000101000;
        10'd170   : cube_lut_2  = 14'b11010000101010;
        10'd171   : cube_lut_2  = 14'b11010000101100;
        10'd172   : cube_lut_2  = 14'b11010000101110;
        10'd173   : cube_lut_2  = 14'b11010000110000;
        10'd174   : cube_lut_2  = 14'b11010000110010;
        10'd175   : cube_lut_2  = 14'b11010000110100;
        10'd176   : cube_lut_2  = 14'b11010000110110;
        10'd177   : cube_lut_2  = 14'b11010000111000;
        10'd178   : cube_lut_2  = 14'b11010000111010;
        10'd179   : cube_lut_2  = 14'b11010000111100;
        10'd180   : cube_lut_2  = 14'b11010000111110;
        10'd181   : cube_lut_2  = 14'b11010001000000;
        10'd182   : cube_lut_2  = 14'b11010001000010;
        10'd183   : cube_lut_2  = 14'b11010001000100;
        10'd184   : cube_lut_2  = 14'b11010001000110;
        10'd185   : cube_lut_2  = 14'b11010001001000;
        10'd186   : cube_lut_2  = 14'b11010001001010;
        10'd187   : cube_lut_2  = 14'b11010001001100;
        10'd188   : cube_lut_2  = 14'b11010001001110;
        10'd189   : cube_lut_2  = 14'b11010001010000;
        10'd190   : cube_lut_2  = 14'b11010001010010;
        10'd191   : cube_lut_2  = 14'b11010001010100;
        10'd192   : cube_lut_2  = 14'b11010001010110;
        10'd193   : cube_lut_2  = 14'b11010001011000;
        10'd194   : cube_lut_2  = 14'b11010001011010;
        10'd195   : cube_lut_2  = 14'b11010001011100;
        10'd196   : cube_lut_2  = 14'b11010001011110;
        10'd197   : cube_lut_2  = 14'b11010001100000;
        10'd198   : cube_lut_2  = 14'b11010001100010;
        10'd199   : cube_lut_2  = 14'b11010001100100;
        10'd200   : cube_lut_2  = 14'b11010001100110;
        10'd201   : cube_lut_2  = 14'b11010001101000;
        10'd202   : cube_lut_2  = 14'b11010001101010;
        10'd203   : cube_lut_2  = 14'b11010001101100;
        10'd204   : cube_lut_2  = 14'b11010001101110;
        10'd205   : cube_lut_2  = 14'b11010001110000;
        10'd206   : cube_lut_2  = 14'b11010001110010;
        10'd207   : cube_lut_2  = 14'b11010001110100;
        10'd208   : cube_lut_2  = 14'b11010001110110;
        10'd209   : cube_lut_2  = 14'b11010001111000;
        10'd210   : cube_lut_2  = 14'b11010001111010;
        10'd211   : cube_lut_2  = 14'b11010001111100;
        10'd212   : cube_lut_2  = 14'b11010001111110;
        10'd213   : cube_lut_2  = 14'b11010010000000;
        10'd214   : cube_lut_2  = 14'b11010010000010;
        10'd215   : cube_lut_2  = 14'b11010010000011;
        10'd216   : cube_lut_2  = 14'b11010010000101;
        10'd217   : cube_lut_2  = 14'b11010010000111;
        10'd218   : cube_lut_2  = 14'b11010010001001;
        10'd219   : cube_lut_2  = 14'b11010010001011;
        10'd220   : cube_lut_2  = 14'b11010010001101;
        10'd221   : cube_lut_2  = 14'b11010010001111;
        10'd222   : cube_lut_2  = 14'b11010010010001;
        10'd223   : cube_lut_2  = 14'b11010010010011;
        10'd224   : cube_lut_2  = 14'b11010010010101;
        10'd225   : cube_lut_2  = 14'b11010010010111;
        10'd226   : cube_lut_2  = 14'b11010010011001;
        10'd227   : cube_lut_2  = 14'b11010010011011;
        10'd228   : cube_lut_2  = 14'b11010010011101;
        10'd229   : cube_lut_2  = 14'b11010010011111;
        10'd230   : cube_lut_2  = 14'b11010010100001;
        10'd231   : cube_lut_2  = 14'b11010010100011;
        10'd232   : cube_lut_2  = 14'b11010010100101;
        10'd233   : cube_lut_2  = 14'b11010010100111;
        10'd234   : cube_lut_2  = 14'b11010010101001;
        10'd235   : cube_lut_2  = 14'b11010010101011;
        10'd236   : cube_lut_2  = 14'b11010010101101;
        10'd237   : cube_lut_2  = 14'b11010010101111;
        10'd238   : cube_lut_2  = 14'b11010010110001;
        10'd239   : cube_lut_2  = 14'b11010010110011;
        10'd240   : cube_lut_2  = 14'b11010010110101;
        10'd241   : cube_lut_2  = 14'b11010010110111;
        10'd242   : cube_lut_2  = 14'b11010010111001;
        10'd243   : cube_lut_2  = 14'b11010010111011;
        10'd244   : cube_lut_2  = 14'b11010010111101;
        10'd245   : cube_lut_2  = 14'b11010010111111;
        10'd246   : cube_lut_2  = 14'b11010011000001;
        10'd247   : cube_lut_2  = 14'b11010011000011;
        10'd248   : cube_lut_2  = 14'b11010011000101;
        10'd249   : cube_lut_2  = 14'b11010011000110;
        10'd250   : cube_lut_2  = 14'b11010011001000;
        10'd251   : cube_lut_2  = 14'b11010011001010;
        10'd252   : cube_lut_2  = 14'b11010011001100;
        10'd253   : cube_lut_2  = 14'b11010011001110;
        10'd254   : cube_lut_2  = 14'b11010011010000;
        10'd255   : cube_lut_2  = 14'b11010011010010;
        10'd256   : cube_lut_2  = 14'b11010011010100;
        10'd257   : cube_lut_2  = 14'b11010011010110;
        10'd258   : cube_lut_2  = 14'b11010011011000;
        10'd259   : cube_lut_2  = 14'b11010011011010;
        10'd260   : cube_lut_2  = 14'b11010011011100;
        10'd261   : cube_lut_2  = 14'b11010011011110;
        10'd262   : cube_lut_2  = 14'b11010011100000;
        10'd263   : cube_lut_2  = 14'b11010011100010;
        10'd264   : cube_lut_2  = 14'b11010011100100;
        10'd265   : cube_lut_2  = 14'b11010011100110;
        10'd266   : cube_lut_2  = 14'b11010011101000;
        10'd267   : cube_lut_2  = 14'b11010011101010;
        10'd268   : cube_lut_2  = 14'b11010011101100;
        10'd269   : cube_lut_2  = 14'b11010011101110;
        10'd270   : cube_lut_2  = 14'b11010011110000;
        10'd271   : cube_lut_2  = 14'b11010011110001;
        10'd272   : cube_lut_2  = 14'b11010011110011;
        10'd273   : cube_lut_2  = 14'b11010011110101;
        10'd274   : cube_lut_2  = 14'b11010011110111;
        10'd275   : cube_lut_2  = 14'b11010011111001;
        10'd276   : cube_lut_2  = 14'b11010011111011;
        10'd277   : cube_lut_2  = 14'b11010011111101;
        10'd278   : cube_lut_2  = 14'b11010011111111;
        10'd279   : cube_lut_2  = 14'b11010100000001;
        10'd280   : cube_lut_2  = 14'b11010100000011;
        10'd281   : cube_lut_2  = 14'b11010100000101;
        10'd282   : cube_lut_2  = 14'b11010100000111;
        10'd283   : cube_lut_2  = 14'b11010100001001;
        10'd284   : cube_lut_2  = 14'b11010100001011;
        10'd285   : cube_lut_2  = 14'b11010100001101;
        10'd286   : cube_lut_2  = 14'b11010100001111;
        10'd287   : cube_lut_2  = 14'b11010100010001;
        10'd288   : cube_lut_2  = 14'b11010100010011;
        10'd289   : cube_lut_2  = 14'b11010100010100;
        10'd290   : cube_lut_2  = 14'b11010100010110;
        10'd291   : cube_lut_2  = 14'b11010100011000;
        10'd292   : cube_lut_2  = 14'b11010100011010;
        10'd293   : cube_lut_2  = 14'b11010100011100;
        10'd294   : cube_lut_2  = 14'b11010100011110;
        10'd295   : cube_lut_2  = 14'b11010100100000;
        10'd296   : cube_lut_2  = 14'b11010100100010;
        10'd297   : cube_lut_2  = 14'b11010100100100;
        10'd298   : cube_lut_2  = 14'b11010100100110;
        10'd299   : cube_lut_2  = 14'b11010100101000;
        10'd300   : cube_lut_2  = 14'b11010100101010;
        10'd301   : cube_lut_2  = 14'b11010100101100;
        10'd302   : cube_lut_2  = 14'b11010100101110;
        10'd303   : cube_lut_2  = 14'b11010100110000;
        10'd304   : cube_lut_2  = 14'b11010100110001;
        10'd305   : cube_lut_2  = 14'b11010100110011;
        10'd306   : cube_lut_2  = 14'b11010100110101;
        10'd307   : cube_lut_2  = 14'b11010100110111;
        10'd308   : cube_lut_2  = 14'b11010100111001;
        10'd309   : cube_lut_2  = 14'b11010100111011;
        10'd310   : cube_lut_2  = 14'b11010100111101;
        10'd311   : cube_lut_2  = 14'b11010100111111;
        10'd312   : cube_lut_2  = 14'b11010101000001;
        10'd313   : cube_lut_2  = 14'b11010101000011;
        10'd314   : cube_lut_2  = 14'b11010101000101;
        10'd315   : cube_lut_2  = 14'b11010101000111;
        10'd316   : cube_lut_2  = 14'b11010101001001;
        10'd317   : cube_lut_2  = 14'b11010101001011;
        10'd318   : cube_lut_2  = 14'b11010101001100;
        10'd319   : cube_lut_2  = 14'b11010101001110;
        10'd320   : cube_lut_2  = 14'b11010101010000;
        10'd321   : cube_lut_2  = 14'b11010101010010;
        10'd322   : cube_lut_2  = 14'b11010101010100;
        10'd323   : cube_lut_2  = 14'b11010101010110;
        10'd324   : cube_lut_2  = 14'b11010101011000;
        10'd325   : cube_lut_2  = 14'b11010101011010;
        10'd326   : cube_lut_2  = 14'b11010101011100;
        10'd327   : cube_lut_2  = 14'b11010101011110;
        10'd328   : cube_lut_2  = 14'b11010101100000;
        10'd329   : cube_lut_2  = 14'b11010101100010;
        10'd330   : cube_lut_2  = 14'b11010101100011;
        10'd331   : cube_lut_2  = 14'b11010101100101;
        10'd332   : cube_lut_2  = 14'b11010101100111;
        10'd333   : cube_lut_2  = 14'b11010101101001;
        10'd334   : cube_lut_2  = 14'b11010101101011;
        10'd335   : cube_lut_2  = 14'b11010101101101;
        10'd336   : cube_lut_2  = 14'b11010101101111;
        10'd337   : cube_lut_2  = 14'b11010101110001;
        10'd338   : cube_lut_2  = 14'b11010101110011;
        10'd339   : cube_lut_2  = 14'b11010101110101;
        10'd340   : cube_lut_2  = 14'b11010101110111;
        10'd341   : cube_lut_2  = 14'b11010101111001;
        10'd342   : cube_lut_2  = 14'b11010101111010;
        10'd343   : cube_lut_2  = 14'b11010101111100;
        10'd344   : cube_lut_2  = 14'b11010101111110;
        10'd345   : cube_lut_2  = 14'b11010110000000;
        10'd346   : cube_lut_2  = 14'b11010110000010;
        10'd347   : cube_lut_2  = 14'b11010110000100;
        10'd348   : cube_lut_2  = 14'b11010110000110;
        10'd349   : cube_lut_2  = 14'b11010110001000;
        10'd350   : cube_lut_2  = 14'b11010110001010;
        10'd351   : cube_lut_2  = 14'b11010110001100;
        10'd352   : cube_lut_2  = 14'b11010110001101;
        10'd353   : cube_lut_2  = 14'b11010110001111;
        10'd354   : cube_lut_2  = 14'b11010110010001;
        10'd355   : cube_lut_2  = 14'b11010110010011;
        10'd356   : cube_lut_2  = 14'b11010110010101;
        10'd357   : cube_lut_2  = 14'b11010110010111;
        10'd358   : cube_lut_2  = 14'b11010110011001;
        10'd359   : cube_lut_2  = 14'b11010110011011;
        10'd360   : cube_lut_2  = 14'b11010110011101;
        10'd361   : cube_lut_2  = 14'b11010110011111;
        10'd362   : cube_lut_2  = 14'b11010110100001;
        10'd363   : cube_lut_2  = 14'b11010110100010;
        10'd364   : cube_lut_2  = 14'b11010110100100;
        10'd365   : cube_lut_2  = 14'b11010110100110;
        10'd366   : cube_lut_2  = 14'b11010110101000;
        10'd367   : cube_lut_2  = 14'b11010110101010;
        10'd368   : cube_lut_2  = 14'b11010110101100;
        10'd369   : cube_lut_2  = 14'b11010110101110;
        10'd370   : cube_lut_2  = 14'b11010110110000;
        10'd371   : cube_lut_2  = 14'b11010110110010;
        10'd372   : cube_lut_2  = 14'b11010110110011;
        10'd373   : cube_lut_2  = 14'b11010110110101;
        10'd374   : cube_lut_2  = 14'b11010110110111;
        10'd375   : cube_lut_2  = 14'b11010110111001;
        10'd376   : cube_lut_2  = 14'b11010110111011;
        10'd377   : cube_lut_2  = 14'b11010110111101;
        10'd378   : cube_lut_2  = 14'b11010110111111;
        10'd379   : cube_lut_2  = 14'b11010111000001;
        10'd380   : cube_lut_2  = 14'b11010111000011;
        10'd381   : cube_lut_2  = 14'b11010111000100;
        10'd382   : cube_lut_2  = 14'b11010111000110;
        10'd383   : cube_lut_2  = 14'b11010111001000;
        10'd384   : cube_lut_2  = 14'b11010111001010;
        10'd385   : cube_lut_2  = 14'b11010111001100;
        10'd386   : cube_lut_2  = 14'b11010111001110;
        10'd387   : cube_lut_2  = 14'b11010111010000;
        10'd388   : cube_lut_2  = 14'b11010111010010;
        10'd389   : cube_lut_2  = 14'b11010111010100;
        10'd390   : cube_lut_2  = 14'b11010111010101;
        10'd391   : cube_lut_2  = 14'b11010111010111;
        10'd392   : cube_lut_2  = 14'b11010111011001;
        10'd393   : cube_lut_2  = 14'b11010111011011;
        10'd394   : cube_lut_2  = 14'b11010111011101;
        10'd395   : cube_lut_2  = 14'b11010111011111;
        10'd396   : cube_lut_2  = 14'b11010111100001;
        10'd397   : cube_lut_2  = 14'b11010111100011;
        10'd398   : cube_lut_2  = 14'b11010111100101;
        10'd399   : cube_lut_2  = 14'b11010111100110;
        10'd400   : cube_lut_2  = 14'b11010111101000;
        10'd401   : cube_lut_2  = 14'b11010111101010;
        10'd402   : cube_lut_2  = 14'b11010111101100;
        10'd403   : cube_lut_2  = 14'b11010111101110;
        10'd404   : cube_lut_2  = 14'b11010111110000;
        10'd405   : cube_lut_2  = 14'b11010111110010;
        10'd406   : cube_lut_2  = 14'b11010111110100;
        10'd407   : cube_lut_2  = 14'b11010111110101;
        10'd408   : cube_lut_2  = 14'b11010111110111;
        10'd409   : cube_lut_2  = 14'b11010111111001;
        10'd410   : cube_lut_2  = 14'b11010111111011;
        10'd411   : cube_lut_2  = 14'b11010111111101;
        10'd412   : cube_lut_2  = 14'b11010111111111;
        10'd413   : cube_lut_2  = 14'b11011000000001;
        10'd414   : cube_lut_2  = 14'b11011000000011;
        10'd415   : cube_lut_2  = 14'b11011000000100;
        10'd416   : cube_lut_2  = 14'b11011000000110;
        10'd417   : cube_lut_2  = 14'b11011000001000;
        10'd418   : cube_lut_2  = 14'b11011000001010;
        10'd419   : cube_lut_2  = 14'b11011000001100;
        10'd420   : cube_lut_2  = 14'b11011000001110;
        10'd421   : cube_lut_2  = 14'b11011000010000;
        10'd422   : cube_lut_2  = 14'b11011000010010;
        10'd423   : cube_lut_2  = 14'b11011000010011;
        10'd424   : cube_lut_2  = 14'b11011000010101;
        10'd425   : cube_lut_2  = 14'b11011000010111;
        10'd426   : cube_lut_2  = 14'b11011000011001;
        10'd427   : cube_lut_2  = 14'b11011000011011;
        10'd428   : cube_lut_2  = 14'b11011000011101;
        10'd429   : cube_lut_2  = 14'b11011000011111;
        10'd430   : cube_lut_2  = 14'b11011000100000;
        10'd431   : cube_lut_2  = 14'b11011000100010;
        10'd432   : cube_lut_2  = 14'b11011000100100;
        10'd433   : cube_lut_2  = 14'b11011000100110;
        10'd434   : cube_lut_2  = 14'b11011000101000;
        10'd435   : cube_lut_2  = 14'b11011000101010;
        10'd436   : cube_lut_2  = 14'b11011000101100;
        10'd437   : cube_lut_2  = 14'b11011000101101;
        10'd438   : cube_lut_2  = 14'b11011000101111;
        10'd439   : cube_lut_2  = 14'b11011000110001;
        10'd440   : cube_lut_2  = 14'b11011000110011;
        10'd441   : cube_lut_2  = 14'b11011000110101;
        10'd442   : cube_lut_2  = 14'b11011000110111;
        10'd443   : cube_lut_2  = 14'b11011000111001;
        10'd444   : cube_lut_2  = 14'b11011000111010;
        10'd445   : cube_lut_2  = 14'b11011000111100;
        10'd446   : cube_lut_2  = 14'b11011000111110;
        10'd447   : cube_lut_2  = 14'b11011001000000;
        10'd448   : cube_lut_2  = 14'b11011001000010;
        10'd449   : cube_lut_2  = 14'b11011001000100;
        10'd450   : cube_lut_2  = 14'b11011001000110;
        10'd451   : cube_lut_2  = 14'b11011001000111;
        10'd452   : cube_lut_2  = 14'b11011001001001;
        10'd453   : cube_lut_2  = 14'b11011001001011;
        10'd454   : cube_lut_2  = 14'b11011001001101;
        10'd455   : cube_lut_2  = 14'b11011001001111;
        10'd456   : cube_lut_2  = 14'b11011001010001;
        10'd457   : cube_lut_2  = 14'b11011001010011;
        10'd458   : cube_lut_2  = 14'b11011001010100;
        10'd459   : cube_lut_2  = 14'b11011001010110;
        10'd460   : cube_lut_2  = 14'b11011001011000;
        10'd461   : cube_lut_2  = 14'b11011001011010;
        10'd462   : cube_lut_2  = 14'b11011001011100;
        10'd463   : cube_lut_2  = 14'b11011001011110;
        10'd464   : cube_lut_2  = 14'b11011001100000;
        10'd465   : cube_lut_2  = 14'b11011001100001;
        10'd466   : cube_lut_2  = 14'b11011001100011;
        10'd467   : cube_lut_2  = 14'b11011001100101;
        10'd468   : cube_lut_2  = 14'b11011001100111;
        10'd469   : cube_lut_2  = 14'b11011001101001;
        10'd470   : cube_lut_2  = 14'b11011001101011;
        10'd471   : cube_lut_2  = 14'b11011001101100;
        10'd472   : cube_lut_2  = 14'b11011001101110;
        10'd473   : cube_lut_2  = 14'b11011001110000;
        10'd474   : cube_lut_2  = 14'b11011001110010;
        10'd475   : cube_lut_2  = 14'b11011001110100;
        10'd476   : cube_lut_2  = 14'b11011001110110;
        10'd477   : cube_lut_2  = 14'b11011001110111;
        10'd478   : cube_lut_2  = 14'b11011001111001;
        10'd479   : cube_lut_2  = 14'b11011001111011;
        10'd480   : cube_lut_2  = 14'b11011001111101;
        10'd481   : cube_lut_2  = 14'b11011001111111;
        10'd482   : cube_lut_2  = 14'b11011010000001;
        10'd483   : cube_lut_2  = 14'b11011010000011;
        10'd484   : cube_lut_2  = 14'b11011010000100;
        10'd485   : cube_lut_2  = 14'b11011010000110;
        10'd486   : cube_lut_2  = 14'b11011010001000;
        10'd487   : cube_lut_2  = 14'b11011010001010;
        10'd488   : cube_lut_2  = 14'b11011010001100;
        10'd489   : cube_lut_2  = 14'b11011010001110;
        10'd490   : cube_lut_2  = 14'b11011010001111;
        10'd491   : cube_lut_2  = 14'b11011010010001;
        10'd492   : cube_lut_2  = 14'b11011010010011;
        10'd493   : cube_lut_2  = 14'b11011010010101;
        10'd494   : cube_lut_2  = 14'b11011010010111;
        10'd495   : cube_lut_2  = 14'b11011010011001;
        10'd496   : cube_lut_2  = 14'b11011010011010;
        10'd497   : cube_lut_2  = 14'b11011010011100;
        10'd498   : cube_lut_2  = 14'b11011010011110;
        10'd499   : cube_lut_2  = 14'b11011010100000;
        10'd500   : cube_lut_2  = 14'b11011010100010;
        10'd501   : cube_lut_2  = 14'b11011010100100;
        10'd502   : cube_lut_2  = 14'b11011010100101;
        10'd503   : cube_lut_2  = 14'b11011010100111;
        10'd504   : cube_lut_2  = 14'b11011010101001;
        10'd505   : cube_lut_2  = 14'b11011010101011;
        10'd506   : cube_lut_2  = 14'b11011010101101;
        10'd507   : cube_lut_2  = 14'b11011010101110;
        10'd508   : cube_lut_2  = 14'b11011010110000;
        10'd509   : cube_lut_2  = 14'b11011010110010;
        10'd510   : cube_lut_2  = 14'b11011010110100;
        10'd511   : cube_lut_2  = 14'b11011010110110;
        10'd512   : cube_lut_2  = 14'b11011010111000;
        10'd513   : cube_lut_2  = 14'b11011010111001;
        10'd514   : cube_lut_2  = 14'b11011010111011;
        10'd515   : cube_lut_2  = 14'b11011010111101;
        10'd516   : cube_lut_2  = 14'b11011010111111;
        10'd517   : cube_lut_2  = 14'b11011011000001;
        10'd518   : cube_lut_2  = 14'b11011011000011;
        10'd519   : cube_lut_2  = 14'b11011011000100;
        10'd520   : cube_lut_2  = 14'b11011011000110;
        10'd521   : cube_lut_2  = 14'b11011011001000;
        10'd522   : cube_lut_2  = 14'b11011011001010;
        10'd523   : cube_lut_2  = 14'b11011011001100;
        10'd524   : cube_lut_2  = 14'b11011011001101;
        10'd525   : cube_lut_2  = 14'b11011011001111;
        10'd526   : cube_lut_2  = 14'b11011011010001;
        10'd527   : cube_lut_2  = 14'b11011011010011;
        10'd528   : cube_lut_2  = 14'b11011011010101;
        10'd529   : cube_lut_2  = 14'b11011011010111;
        10'd530   : cube_lut_2  = 14'b11011011011000;
        10'd531   : cube_lut_2  = 14'b11011011011010;
        10'd532   : cube_lut_2  = 14'b11011011011100;
        10'd533   : cube_lut_2  = 14'b11011011011110;
        10'd534   : cube_lut_2  = 14'b11011011100000;
        10'd535   : cube_lut_2  = 14'b11011011100001;
        10'd536   : cube_lut_2  = 14'b11011011100011;
        10'd537   : cube_lut_2  = 14'b11011011100101;
        10'd538   : cube_lut_2  = 14'b11011011100111;
        10'd539   : cube_lut_2  = 14'b11011011101001;
        10'd540   : cube_lut_2  = 14'b11011011101011;
        10'd541   : cube_lut_2  = 14'b11011011101100;
        10'd542   : cube_lut_2  = 14'b11011011101110;
        10'd543   : cube_lut_2  = 14'b11011011110000;
        10'd544   : cube_lut_2  = 14'b11011011110010;
        10'd545   : cube_lut_2  = 14'b11011011110100;
        10'd546   : cube_lut_2  = 14'b11011011110101;
        10'd547   : cube_lut_2  = 14'b11011011110111;
        10'd548   : cube_lut_2  = 14'b11011011111001;
        10'd549   : cube_lut_2  = 14'b11011011111011;
        10'd550   : cube_lut_2  = 14'b11011011111101;
        10'd551   : cube_lut_2  = 14'b11011011111110;
        10'd552   : cube_lut_2  = 14'b11011100000000;
        10'd553   : cube_lut_2  = 14'b11011100000010;
        10'd554   : cube_lut_2  = 14'b11011100000100;
        10'd555   : cube_lut_2  = 14'b11011100000110;
        10'd556   : cube_lut_2  = 14'b11011100000111;
        10'd557   : cube_lut_2  = 14'b11011100001001;
        10'd558   : cube_lut_2  = 14'b11011100001011;
        10'd559   : cube_lut_2  = 14'b11011100001101;
        10'd560   : cube_lut_2  = 14'b11011100001111;
        10'd561   : cube_lut_2  = 14'b11011100010000;
        10'd562   : cube_lut_2  = 14'b11011100010010;
        10'd563   : cube_lut_2  = 14'b11011100010100;
        10'd564   : cube_lut_2  = 14'b11011100010110;
        10'd565   : cube_lut_2  = 14'b11011100011000;
        10'd566   : cube_lut_2  = 14'b11011100011001;
        10'd567   : cube_lut_2  = 14'b11011100011011;
        10'd568   : cube_lut_2  = 14'b11011100011101;
        10'd569   : cube_lut_2  = 14'b11011100011111;
        10'd570   : cube_lut_2  = 14'b11011100100001;
        10'd571   : cube_lut_2  = 14'b11011100100010;
        10'd572   : cube_lut_2  = 14'b11011100100100;
        10'd573   : cube_lut_2  = 14'b11011100100110;
        10'd574   : cube_lut_2  = 14'b11011100101000;
        10'd575   : cube_lut_2  = 14'b11011100101010;
        10'd576   : cube_lut_2  = 14'b11011100101011;
        10'd577   : cube_lut_2  = 14'b11011100101101;
        10'd578   : cube_lut_2  = 14'b11011100101111;
        10'd579   : cube_lut_2  = 14'b11011100110001;
        10'd580   : cube_lut_2  = 14'b11011100110011;
        10'd581   : cube_lut_2  = 14'b11011100110100;
        10'd582   : cube_lut_2  = 14'b11011100110110;
        10'd583   : cube_lut_2  = 14'b11011100111000;
        10'd584   : cube_lut_2  = 14'b11011100111010;
        10'd585   : cube_lut_2  = 14'b11011100111100;
        10'd586   : cube_lut_2  = 14'b11011100111101;
        10'd587   : cube_lut_2  = 14'b11011100111111;
        10'd588   : cube_lut_2  = 14'b11011101000001;
        10'd589   : cube_lut_2  = 14'b11011101000011;
        10'd590   : cube_lut_2  = 14'b11011101000100;
        10'd591   : cube_lut_2  = 14'b11011101000110;
        10'd592   : cube_lut_2  = 14'b11011101001000;
        10'd593   : cube_lut_2  = 14'b11011101001010;
        10'd594   : cube_lut_2  = 14'b11011101001100;
        10'd595   : cube_lut_2  = 14'b11011101001101;
        10'd596   : cube_lut_2  = 14'b11011101001111;
        10'd597   : cube_lut_2  = 14'b11011101010001;
        10'd598   : cube_lut_2  = 14'b11011101010011;
        10'd599   : cube_lut_2  = 14'b11011101010101;
        10'd600   : cube_lut_2  = 14'b11011101010110;
        10'd601   : cube_lut_2  = 14'b11011101011000;
        10'd602   : cube_lut_2  = 14'b11011101011010;
        10'd603   : cube_lut_2  = 14'b11011101011100;
        10'd604   : cube_lut_2  = 14'b11011101011101;
        10'd605   : cube_lut_2  = 14'b11011101011111;
        10'd606   : cube_lut_2  = 14'b11011101100001;
        10'd607   : cube_lut_2  = 14'b11011101100011;
        10'd608   : cube_lut_2  = 14'b11011101100101;
        10'd609   : cube_lut_2  = 14'b11011101100110;
        10'd610   : cube_lut_2  = 14'b11011101101000;
        10'd611   : cube_lut_2  = 14'b11011101101010;
        10'd612   : cube_lut_2  = 14'b11011101101100;
        10'd613   : cube_lut_2  = 14'b11011101101101;
        10'd614   : cube_lut_2  = 14'b11011101101111;
        10'd615   : cube_lut_2  = 14'b11011101110001;
        10'd616   : cube_lut_2  = 14'b11011101110011;
        10'd617   : cube_lut_2  = 14'b11011101110101;
        10'd618   : cube_lut_2  = 14'b11011101110110;
        10'd619   : cube_lut_2  = 14'b11011101111000;
        10'd620   : cube_lut_2  = 14'b11011101111010;
        10'd621   : cube_lut_2  = 14'b11011101111100;
        10'd622   : cube_lut_2  = 14'b11011101111101;
        10'd623   : cube_lut_2  = 14'b11011101111111;
        10'd624   : cube_lut_2  = 14'b11011110000001;
        10'd625   : cube_lut_2  = 14'b11011110000011;
        10'd626   : cube_lut_2  = 14'b11011110000101;
        10'd627   : cube_lut_2  = 14'b11011110000110;
        10'd628   : cube_lut_2  = 14'b11011110001000;
        10'd629   : cube_lut_2  = 14'b11011110001010;
        10'd630   : cube_lut_2  = 14'b11011110001100;
        10'd631   : cube_lut_2  = 14'b11011110001101;
        10'd632   : cube_lut_2  = 14'b11011110001111;
        10'd633   : cube_lut_2  = 14'b11011110010001;
        10'd634   : cube_lut_2  = 14'b11011110010011;
        10'd635   : cube_lut_2  = 14'b11011110010100;
        10'd636   : cube_lut_2  = 14'b11011110010110;
        10'd637   : cube_lut_2  = 14'b11011110011000;
        10'd638   : cube_lut_2  = 14'b11011110011010;
        10'd639   : cube_lut_2  = 14'b11011110011100;
        10'd640   : cube_lut_2  = 14'b11011110011101;
        10'd641   : cube_lut_2  = 14'b11011110011111;
        10'd642   : cube_lut_2  = 14'b11011110100001;
        10'd643   : cube_lut_2  = 14'b11011110100011;
        10'd644   : cube_lut_2  = 14'b11011110100100;
        10'd645   : cube_lut_2  = 14'b11011110100110;
        10'd646   : cube_lut_2  = 14'b11011110101000;
        10'd647   : cube_lut_2  = 14'b11011110101010;
        10'd648   : cube_lut_2  = 14'b11011110101011;
        10'd649   : cube_lut_2  = 14'b11011110101101;
        10'd650   : cube_lut_2  = 14'b11011110101111;
        10'd651   : cube_lut_2  = 14'b11011110110001;
        10'd652   : cube_lut_2  = 14'b11011110110010;
        10'd653   : cube_lut_2  = 14'b11011110110100;
        10'd654   : cube_lut_2  = 14'b11011110110110;
        10'd655   : cube_lut_2  = 14'b11011110111000;
        10'd656   : cube_lut_2  = 14'b11011110111001;
        10'd657   : cube_lut_2  = 14'b11011110111011;
        10'd658   : cube_lut_2  = 14'b11011110111101;
        10'd659   : cube_lut_2  = 14'b11011110111111;
        10'd660   : cube_lut_2  = 14'b11011111000001;
        10'd661   : cube_lut_2  = 14'b11011111000010;
        10'd662   : cube_lut_2  = 14'b11011111000100;
        10'd663   : cube_lut_2  = 14'b11011111000110;
        10'd664   : cube_lut_2  = 14'b11011111001000;
        10'd665   : cube_lut_2  = 14'b11011111001001;
        10'd666   : cube_lut_2  = 14'b11011111001011;
        10'd667   : cube_lut_2  = 14'b11011111001101;
        10'd668   : cube_lut_2  = 14'b11011111001111;
        10'd669   : cube_lut_2  = 14'b11011111010000;
        10'd670   : cube_lut_2  = 14'b11011111010010;
        10'd671   : cube_lut_2  = 14'b11011111010100;
        10'd672   : cube_lut_2  = 14'b11011111010110;
        10'd673   : cube_lut_2  = 14'b11011111010111;
        10'd674   : cube_lut_2  = 14'b11011111011001;
        10'd675   : cube_lut_2  = 14'b11011111011011;
        10'd676   : cube_lut_2  = 14'b11011111011101;
        10'd677   : cube_lut_2  = 14'b11011111011110;
        10'd678   : cube_lut_2  = 14'b11011111100000;
        10'd679   : cube_lut_2  = 14'b11011111100010;
        10'd680   : cube_lut_2  = 14'b11011111100100;
        10'd681   : cube_lut_2  = 14'b11011111100101;
        10'd682   : cube_lut_2  = 14'b11011111100111;
        10'd683   : cube_lut_2  = 14'b11011111101001;
        10'd684   : cube_lut_2  = 14'b11011111101011;
        10'd685   : cube_lut_2  = 14'b11011111101100;
        10'd686   : cube_lut_2  = 14'b11011111101110;
        10'd687   : cube_lut_2  = 14'b11011111110000;
        10'd688   : cube_lut_2  = 14'b11011111110010;
        10'd689   : cube_lut_2  = 14'b11011111110011;
        10'd690   : cube_lut_2  = 14'b11011111110101;
        10'd691   : cube_lut_2  = 14'b11011111110111;
        10'd692   : cube_lut_2  = 14'b11011111111001;
        10'd693   : cube_lut_2  = 14'b11011111111010;
        10'd694   : cube_lut_2  = 14'b11011111111100;
        10'd695   : cube_lut_2  = 14'b11011111111110;
        10'd696   : cube_lut_2  = 14'b11100000000000;
        10'd697   : cube_lut_2  = 14'b11100000000001;
        10'd698   : cube_lut_2  = 14'b11100000000011;
        10'd699   : cube_lut_2  = 14'b11100000000101;
        10'd700   : cube_lut_2  = 14'b11100000000110;
        10'd701   : cube_lut_2  = 14'b11100000001000;
        10'd702   : cube_lut_2  = 14'b11100000001010;
        10'd703   : cube_lut_2  = 14'b11100000001100;
        10'd704   : cube_lut_2  = 14'b11100000001101;
        10'd705   : cube_lut_2  = 14'b11100000001111;
        10'd706   : cube_lut_2  = 14'b11100000010001;
        10'd707   : cube_lut_2  = 14'b11100000010011;
        10'd708   : cube_lut_2  = 14'b11100000010100;
        10'd709   : cube_lut_2  = 14'b11100000010110;
        10'd710   : cube_lut_2  = 14'b11100000011000;
        10'd711   : cube_lut_2  = 14'b11100000011010;
        10'd712   : cube_lut_2  = 14'b11100000011011;
        10'd713   : cube_lut_2  = 14'b11100000011101;
        10'd714   : cube_lut_2  = 14'b11100000011111;
        10'd715   : cube_lut_2  = 14'b11100000100001;
        10'd716   : cube_lut_2  = 14'b11100000100010;
        10'd717   : cube_lut_2  = 14'b11100000100100;
        10'd718   : cube_lut_2  = 14'b11100000100110;
        10'd719   : cube_lut_2  = 14'b11100000100111;
        10'd720   : cube_lut_2  = 14'b11100000101001;
        10'd721   : cube_lut_2  = 14'b11100000101011;
        10'd722   : cube_lut_2  = 14'b11100000101101;
        10'd723   : cube_lut_2  = 14'b11100000101110;
        10'd724   : cube_lut_2  = 14'b11100000110000;
        10'd725   : cube_lut_2  = 14'b11100000110010;
        10'd726   : cube_lut_2  = 14'b11100000110100;
        10'd727   : cube_lut_2  = 14'b11100000110101;
        10'd728   : cube_lut_2  = 14'b11100000110111;
        10'd729   : cube_lut_2  = 14'b11100000111001;
        10'd730   : cube_lut_2  = 14'b11100000111010;
        10'd731   : cube_lut_2  = 14'b11100000111100;
        10'd732   : cube_lut_2  = 14'b11100000111110;
        10'd733   : cube_lut_2  = 14'b11100001000000;
        10'd734   : cube_lut_2  = 14'b11100001000001;
        10'd735   : cube_lut_2  = 14'b11100001000011;
        10'd736   : cube_lut_2  = 14'b11100001000101;
        10'd737   : cube_lut_2  = 14'b11100001000111;
        10'd738   : cube_lut_2  = 14'b11100001001000;
        10'd739   : cube_lut_2  = 14'b11100001001010;
        10'd740   : cube_lut_2  = 14'b11100001001100;
        10'd741   : cube_lut_2  = 14'b11100001001101;
        10'd742   : cube_lut_2  = 14'b11100001001111;
        10'd743   : cube_lut_2  = 14'b11100001010001;
        10'd744   : cube_lut_2  = 14'b11100001010011;
        10'd745   : cube_lut_2  = 14'b11100001010100;
        10'd746   : cube_lut_2  = 14'b11100001010110;
        10'd747   : cube_lut_2  = 14'b11100001011000;
        10'd748   : cube_lut_2  = 14'b11100001011001;
        10'd749   : cube_lut_2  = 14'b11100001011011;
        10'd750   : cube_lut_2  = 14'b11100001011101;
        10'd751   : cube_lut_2  = 14'b11100001011111;
        10'd752   : cube_lut_2  = 14'b11100001100000;
        10'd753   : cube_lut_2  = 14'b11100001100010;
        10'd754   : cube_lut_2  = 14'b11100001100100;
        10'd755   : cube_lut_2  = 14'b11100001100110;
        10'd756   : cube_lut_2  = 14'b11100001100111;
        10'd757   : cube_lut_2  = 14'b11100001101001;
        10'd758   : cube_lut_2  = 14'b11100001101011;
        10'd759   : cube_lut_2  = 14'b11100001101100;
        10'd760   : cube_lut_2  = 14'b11100001101110;
        10'd761   : cube_lut_2  = 14'b11100001110000;
        10'd762   : cube_lut_2  = 14'b11100001110010;
        10'd763   : cube_lut_2  = 14'b11100001110011;
        10'd764   : cube_lut_2  = 14'b11100001110101;
        10'd765   : cube_lut_2  = 14'b11100001110111;
        10'd766   : cube_lut_2  = 14'b11100001111000;
        10'd767   : cube_lut_2  = 14'b11100001111010;
        10'd768   : cube_lut_2  = 14'b11100001111100;
        10'd769   : cube_lut_2  = 14'b11100001111110;
        10'd770   : cube_lut_2  = 14'b11100001111111;
        10'd771   : cube_lut_2  = 14'b11100010000001;
        10'd772   : cube_lut_2  = 14'b11100010000011;
        10'd773   : cube_lut_2  = 14'b11100010000100;
        10'd774   : cube_lut_2  = 14'b11100010000110;
        10'd775   : cube_lut_2  = 14'b11100010001000;
        10'd776   : cube_lut_2  = 14'b11100010001001;
        10'd777   : cube_lut_2  = 14'b11100010001011;
        10'd778   : cube_lut_2  = 14'b11100010001101;
        10'd779   : cube_lut_2  = 14'b11100010001111;
        10'd780   : cube_lut_2  = 14'b11100010010000;
        10'd781   : cube_lut_2  = 14'b11100010010010;
        10'd782   : cube_lut_2  = 14'b11100010010100;
        10'd783   : cube_lut_2  = 14'b11100010010101;
        10'd784   : cube_lut_2  = 14'b11100010010111;
        10'd785   : cube_lut_2  = 14'b11100010011001;
        10'd786   : cube_lut_2  = 14'b11100010011011;
        10'd787   : cube_lut_2  = 14'b11100010011100;
        10'd788   : cube_lut_2  = 14'b11100010011110;
        10'd789   : cube_lut_2  = 14'b11100010100000;
        10'd790   : cube_lut_2  = 14'b11100010100001;
        10'd791   : cube_lut_2  = 14'b11100010100011;
        10'd792   : cube_lut_2  = 14'b11100010100101;
        10'd793   : cube_lut_2  = 14'b11100010100110;
        10'd794   : cube_lut_2  = 14'b11100010101000;
        10'd795   : cube_lut_2  = 14'b11100010101010;
        10'd796   : cube_lut_2  = 14'b11100010101100;
        10'd797   : cube_lut_2  = 14'b11100010101101;
        10'd798   : cube_lut_2  = 14'b11100010101111;
        10'd799   : cube_lut_2  = 14'b11100010110001;
        10'd800   : cube_lut_2  = 14'b11100010110010;
        10'd801   : cube_lut_2  = 14'b11100010110100;
        10'd802   : cube_lut_2  = 14'b11100010110110;
        10'd803   : cube_lut_2  = 14'b11100010110111;
        10'd804   : cube_lut_2  = 14'b11100010111001;
        10'd805   : cube_lut_2  = 14'b11100010111011;
        10'd806   : cube_lut_2  = 14'b11100010111101;
        10'd807   : cube_lut_2  = 14'b11100010111110;
        10'd808   : cube_lut_2  = 14'b11100011000000;
        10'd809   : cube_lut_2  = 14'b11100011000010;
        10'd810   : cube_lut_2  = 14'b11100011000011;
        10'd811   : cube_lut_2  = 14'b11100011000101;
        10'd812   : cube_lut_2  = 14'b11100011000111;
        10'd813   : cube_lut_2  = 14'b11100011001000;
        10'd814   : cube_lut_2  = 14'b11100011001010;
        10'd815   : cube_lut_2  = 14'b11100011001100;
        10'd816   : cube_lut_2  = 14'b11100011001110;
        10'd817   : cube_lut_2  = 14'b11100011001111;
        10'd818   : cube_lut_2  = 14'b11100011010001;
        10'd819   : cube_lut_2  = 14'b11100011010011;
        10'd820   : cube_lut_2  = 14'b11100011010100;
        10'd821   : cube_lut_2  = 14'b11100011010110;
        10'd822   : cube_lut_2  = 14'b11100011011000;
        10'd823   : cube_lut_2  = 14'b11100011011001;
        10'd824   : cube_lut_2  = 14'b11100011011011;
        10'd825   : cube_lut_2  = 14'b11100011011101;
        10'd826   : cube_lut_2  = 14'b11100011011110;
        10'd827   : cube_lut_2  = 14'b11100011100000;
        10'd828   : cube_lut_2  = 14'b11100011100010;
        10'd829   : cube_lut_2  = 14'b11100011100011;
        10'd830   : cube_lut_2  = 14'b11100011100101;
        10'd831   : cube_lut_2  = 14'b11100011100111;
        10'd832   : cube_lut_2  = 14'b11100011101001;
        10'd833   : cube_lut_2  = 14'b11100011101010;
        10'd834   : cube_lut_2  = 14'b11100011101100;
        10'd835   : cube_lut_2  = 14'b11100011101110;
        10'd836   : cube_lut_2  = 14'b11100011101111;
        10'd837   : cube_lut_2  = 14'b11100011110001;
        10'd838   : cube_lut_2  = 14'b11100011110011;
        10'd839   : cube_lut_2  = 14'b11100011110100;
        10'd840   : cube_lut_2  = 14'b11100011110110;
        10'd841   : cube_lut_2  = 14'b11100011111000;
        10'd842   : cube_lut_2  = 14'b11100011111001;
        10'd843   : cube_lut_2  = 14'b11100011111011;
        10'd844   : cube_lut_2  = 14'b11100011111101;
        10'd845   : cube_lut_2  = 14'b11100011111110;
        10'd846   : cube_lut_2  = 14'b11100100000000;
        10'd847   : cube_lut_2  = 14'b11100100000010;
        10'd848   : cube_lut_2  = 14'b11100100000011;
        10'd849   : cube_lut_2  = 14'b11100100000101;
        10'd850   : cube_lut_2  = 14'b11100100000111;
        10'd851   : cube_lut_2  = 14'b11100100001001;
        10'd852   : cube_lut_2  = 14'b11100100001010;
        10'd853   : cube_lut_2  = 14'b11100100001100;
        10'd854   : cube_lut_2  = 14'b11100100001110;
        10'd855   : cube_lut_2  = 14'b11100100001111;
        10'd856   : cube_lut_2  = 14'b11100100010001;
        10'd857   : cube_lut_2  = 14'b11100100010011;
        10'd858   : cube_lut_2  = 14'b11100100010100;
        10'd859   : cube_lut_2  = 14'b11100100010110;
        10'd860   : cube_lut_2  = 14'b11100100011000;
        10'd861   : cube_lut_2  = 14'b11100100011001;
        10'd862   : cube_lut_2  = 14'b11100100011011;
        10'd863   : cube_lut_2  = 14'b11100100011101;
        10'd864   : cube_lut_2  = 14'b11100100011110;
        10'd865   : cube_lut_2  = 14'b11100100100000;
        10'd866   : cube_lut_2  = 14'b11100100100010;
        10'd867   : cube_lut_2  = 14'b11100100100011;
        10'd868   : cube_lut_2  = 14'b11100100100101;
        10'd869   : cube_lut_2  = 14'b11100100100111;
        10'd870   : cube_lut_2  = 14'b11100100101000;
        10'd871   : cube_lut_2  = 14'b11100100101010;
        10'd872   : cube_lut_2  = 14'b11100100101100;
        10'd873   : cube_lut_2  = 14'b11100100101101;
        10'd874   : cube_lut_2  = 14'b11100100101111;
        10'd875   : cube_lut_2  = 14'b11100100110001;
        10'd876   : cube_lut_2  = 14'b11100100110010;
        10'd877   : cube_lut_2  = 14'b11100100110100;
        10'd878   : cube_lut_2  = 14'b11100100110110;
        10'd879   : cube_lut_2  = 14'b11100100110111;
        10'd880   : cube_lut_2  = 14'b11100100111001;
        10'd881   : cube_lut_2  = 14'b11100100111011;
        10'd882   : cube_lut_2  = 14'b11100100111100;
        10'd883   : cube_lut_2  = 14'b11100100111110;
        10'd884   : cube_lut_2  = 14'b11100101000000;
        10'd885   : cube_lut_2  = 14'b11100101000001;
        10'd886   : cube_lut_2  = 14'b11100101000011;
        10'd887   : cube_lut_2  = 14'b11100101000101;
        10'd888   : cube_lut_2  = 14'b11100101000110;
        10'd889   : cube_lut_2  = 14'b11100101001000;
        10'd890   : cube_lut_2  = 14'b11100101001010;
        10'd891   : cube_lut_2  = 14'b11100101001011;
        10'd892   : cube_lut_2  = 14'b11100101001101;
        10'd893   : cube_lut_2  = 14'b11100101001111;
        10'd894   : cube_lut_2  = 14'b11100101010000;
        10'd895   : cube_lut_2  = 14'b11100101010010;
        10'd896   : cube_lut_2  = 14'b11100101010100;
        10'd897   : cube_lut_2  = 14'b11100101010101;
        10'd898   : cube_lut_2  = 14'b11100101010111;
        10'd899   : cube_lut_2  = 14'b11100101011001;
        10'd900   : cube_lut_2  = 14'b11100101011010;
        10'd901   : cube_lut_2  = 14'b11100101011100;
        10'd902   : cube_lut_2  = 14'b11100101011110;
        10'd903   : cube_lut_2  = 14'b11100101011111;
        10'd904   : cube_lut_2  = 14'b11100101100001;
        10'd905   : cube_lut_2  = 14'b11100101100011;
        10'd906   : cube_lut_2  = 14'b11100101100100;
        10'd907   : cube_lut_2  = 14'b11100101100110;
        10'd908   : cube_lut_2  = 14'b11100101101000;
        10'd909   : cube_lut_2  = 14'b11100101101001;
        10'd910   : cube_lut_2  = 14'b11100101101011;
        10'd911   : cube_lut_2  = 14'b11100101101101;
        10'd912   : cube_lut_2  = 14'b11100101101110;
        10'd913   : cube_lut_2  = 14'b11100101110000;
        10'd914   : cube_lut_2  = 14'b11100101110010;
        10'd915   : cube_lut_2  = 14'b11100101110011;
        10'd916   : cube_lut_2  = 14'b11100101110101;
        10'd917   : cube_lut_2  = 14'b11100101110110;
        10'd918   : cube_lut_2  = 14'b11100101111000;
        10'd919   : cube_lut_2  = 14'b11100101111010;
        10'd920   : cube_lut_2  = 14'b11100101111011;
        10'd921   : cube_lut_2  = 14'b11100101111101;
        10'd922   : cube_lut_2  = 14'b11100101111111;
        10'd923   : cube_lut_2  = 14'b11100110000000;
        10'd924   : cube_lut_2  = 14'b11100110000010;
        10'd925   : cube_lut_2  = 14'b11100110000100;
        10'd926   : cube_lut_2  = 14'b11100110000101;
        10'd927   : cube_lut_2  = 14'b11100110000111;
        10'd928   : cube_lut_2  = 14'b11100110001001;
        10'd929   : cube_lut_2  = 14'b11100110001010;
        10'd930   : cube_lut_2  = 14'b11100110001100;
        10'd931   : cube_lut_2  = 14'b11100110001110;
        10'd932   : cube_lut_2  = 14'b11100110001111;
        10'd933   : cube_lut_2  = 14'b11100110010001;
        10'd934   : cube_lut_2  = 14'b11100110010011;
        10'd935   : cube_lut_2  = 14'b11100110010100;
        10'd936   : cube_lut_2  = 14'b11100110010110;
        10'd937   : cube_lut_2  = 14'b11100110010111;
        10'd938   : cube_lut_2  = 14'b11100110011001;
        10'd939   : cube_lut_2  = 14'b11100110011011;
        10'd940   : cube_lut_2  = 14'b11100110011100;
        10'd941   : cube_lut_2  = 14'b11100110011110;
        10'd942   : cube_lut_2  = 14'b11100110100000;
        10'd943   : cube_lut_2  = 14'b11100110100001;
        10'd944   : cube_lut_2  = 14'b11100110100011;
        10'd945   : cube_lut_2  = 14'b11100110100101;
        10'd946   : cube_lut_2  = 14'b11100110100110;
        10'd947   : cube_lut_2  = 14'b11100110101000;
        10'd948   : cube_lut_2  = 14'b11100110101010;
        10'd949   : cube_lut_2  = 14'b11100110101011;
        10'd950   : cube_lut_2  = 14'b11100110101101;
        10'd951   : cube_lut_2  = 14'b11100110101110;
        10'd952   : cube_lut_2  = 14'b11100110110000;
        10'd953   : cube_lut_2  = 14'b11100110110010;
        10'd954   : cube_lut_2  = 14'b11100110110011;
        10'd955   : cube_lut_2  = 14'b11100110110101;
        10'd956   : cube_lut_2  = 14'b11100110110111;
        10'd957   : cube_lut_2  = 14'b11100110111000;
        10'd958   : cube_lut_2  = 14'b11100110111010;
        10'd959   : cube_lut_2  = 14'b11100110111100;
        10'd960   : cube_lut_2  = 14'b11100110111101;
        10'd961   : cube_lut_2  = 14'b11100110111111;
        10'd962   : cube_lut_2  = 14'b11100111000001;
        10'd963   : cube_lut_2  = 14'b11100111000010;
        10'd964   : cube_lut_2  = 14'b11100111000100;
        10'd965   : cube_lut_2  = 14'b11100111000101;
        10'd966   : cube_lut_2  = 14'b11100111000111;
        10'd967   : cube_lut_2  = 14'b11100111001001;
        10'd968   : cube_lut_2  = 14'b11100111001010;
        10'd969   : cube_lut_2  = 14'b11100111001100;
        10'd970   : cube_lut_2  = 14'b11100111001110;
        10'd971   : cube_lut_2  = 14'b11100111001111;
        10'd972   : cube_lut_2  = 14'b11100111010001;
        10'd973   : cube_lut_2  = 14'b11100111010011;
        10'd974   : cube_lut_2  = 14'b11100111010100;
        10'd975   : cube_lut_2  = 14'b11100111010110;
        10'd976   : cube_lut_2  = 14'b11100111010111;
        10'd977   : cube_lut_2  = 14'b11100111011001;
        10'd978   : cube_lut_2  = 14'b11100111011011;
        10'd979   : cube_lut_2  = 14'b11100111011100;
        10'd980   : cube_lut_2  = 14'b11100111011110;
        10'd981   : cube_lut_2  = 14'b11100111100000;
        10'd982   : cube_lut_2  = 14'b11100111100001;
        10'd983   : cube_lut_2  = 14'b11100111100011;
        10'd984   : cube_lut_2  = 14'b11100111100100;
        10'd985   : cube_lut_2  = 14'b11100111100110;
        10'd986   : cube_lut_2  = 14'b11100111101000;
        10'd987   : cube_lut_2  = 14'b11100111101001;
        10'd988   : cube_lut_2  = 14'b11100111101011;
        10'd989   : cube_lut_2  = 14'b11100111101101;
        10'd990   : cube_lut_2  = 14'b11100111101110;
        10'd991   : cube_lut_2  = 14'b11100111110000;
        10'd992   : cube_lut_2  = 14'b11100111110001;
        10'd993   : cube_lut_2  = 14'b11100111110011;
        10'd994   : cube_lut_2  = 14'b11100111110101;
        10'd995   : cube_lut_2  = 14'b11100111110110;
        10'd996   : cube_lut_2  = 14'b11100111111000;
        10'd997   : cube_lut_2  = 14'b11100111111010;
        10'd998   : cube_lut_2  = 14'b11100111111011;
        10'd999   : cube_lut_2  = 14'b11100111111101;
        10'd1000   : cube_lut_2 = 14'b11100111111110;
        10'd1001   : cube_lut_2 = 14'b11101000000000;
        10'd1002   : cube_lut_2 = 14'b11101000000010;
        10'd1003   : cube_lut_2 = 14'b11101000000011;
        10'd1004   : cube_lut_2 = 14'b11101000000101;
        10'd1005   : cube_lut_2 = 14'b11101000000111;
        10'd1006   : cube_lut_2 = 14'b11101000001000;
        10'd1007   : cube_lut_2 = 14'b11101000001010;
        10'd1008   : cube_lut_2 = 14'b11101000001011;
        10'd1009   : cube_lut_2 = 14'b11101000001101;
        10'd1010   : cube_lut_2 = 14'b11101000001111;
        10'd1011   : cube_lut_2 = 14'b11101000010000;
        10'd1012   : cube_lut_2 = 14'b11101000010010;
        10'd1013   : cube_lut_2 = 14'b11101000010100;
        10'd1014   : cube_lut_2 = 14'b11101000010101;
        10'd1015   : cube_lut_2 = 14'b11101000010111;
        10'd1016   : cube_lut_2 = 14'b11101000011000;
        10'd1017   : cube_lut_2 = 14'b11101000011010;
        10'd1018   : cube_lut_2 = 14'b11101000011100;
        10'd1019   : cube_lut_2 = 14'b11101000011101;
        10'd1020   : cube_lut_2 = 14'b11101000011111;
        10'd1021   : cube_lut_2 = 14'b11101000100001;
        10'd1022   : cube_lut_2 = 14'b11101000100010;
        10'd1023   : cube_lut_2 = 14'b11101000100100;
        
    endcase
end

always@* begin
    
    cube_lut_3 = 0;
    
    case(i_data[9:0])
        
        10'd0   : cube_lut_3    = 14'b11101000100101;
        10'd1   : cube_lut_3    = 14'b11101000100111;
        10'd2   : cube_lut_3    = 14'b11101000101001;
        10'd3   : cube_lut_3    = 14'b11101000101010;
        10'd4   : cube_lut_3    = 14'b11101000101100;
        10'd5   : cube_lut_3    = 14'b11101000101101;
        10'd6   : cube_lut_3    = 14'b11101000101111;
        10'd7   : cube_lut_3    = 14'b11101000110001;
        10'd8   : cube_lut_3    = 14'b11101000110010;
        10'd9   : cube_lut_3    = 14'b11101000110100;
        10'd10   : cube_lut_3   = 14'b11101000110101;
        10'd11   : cube_lut_3   = 14'b11101000110111;
        10'd12   : cube_lut_3   = 14'b11101000111001;
        10'd13   : cube_lut_3   = 14'b11101000111010;
        10'd14   : cube_lut_3   = 14'b11101000111100;
        10'd15   : cube_lut_3   = 14'b11101000111110;
        10'd16   : cube_lut_3   = 14'b11101000111111;
        10'd17   : cube_lut_3   = 14'b11101001000001;
        10'd18   : cube_lut_3   = 14'b11101001000010;
        10'd19   : cube_lut_3   = 14'b11101001000100;
        10'd20   : cube_lut_3   = 14'b11101001000110;
        10'd21   : cube_lut_3   = 14'b11101001000111;
        10'd22   : cube_lut_3   = 14'b11101001001001;
        10'd23   : cube_lut_3   = 14'b11101001001010;
        10'd24   : cube_lut_3   = 14'b11101001001100;
        10'd25   : cube_lut_3   = 14'b11101001001110;
        10'd26   : cube_lut_3   = 14'b11101001001111;
        10'd27   : cube_lut_3   = 14'b11101001010001;
        10'd28   : cube_lut_3   = 14'b11101001010010;
        10'd29   : cube_lut_3   = 14'b11101001010100;
        10'd30   : cube_lut_3   = 14'b11101001010110;
        10'd31   : cube_lut_3   = 14'b11101001010111;
        10'd32   : cube_lut_3   = 14'b11101001011001;
        10'd33   : cube_lut_3   = 14'b11101001011010;
        10'd34   : cube_lut_3   = 14'b11101001011100;
        10'd35   : cube_lut_3   = 14'b11101001011110;
        10'd36   : cube_lut_3   = 14'b11101001011111;
        10'd37   : cube_lut_3   = 14'b11101001100001;
        10'd38   : cube_lut_3   = 14'b11101001100010;
        10'd39   : cube_lut_3   = 14'b11101001100100;
        10'd40   : cube_lut_3   = 14'b11101001100110;
        10'd41   : cube_lut_3   = 14'b11101001100111;
        10'd42   : cube_lut_3   = 14'b11101001101001;
        10'd43   : cube_lut_3   = 14'b11101001101010;
        10'd44   : cube_lut_3   = 14'b11101001101100;
        10'd45   : cube_lut_3   = 14'b11101001101110;
        10'd46   : cube_lut_3   = 14'b11101001101111;
        10'd47   : cube_lut_3   = 14'b11101001110001;
        10'd48   : cube_lut_3   = 14'b11101001110010;
        10'd49   : cube_lut_3   = 14'b11101001110100;
        10'd50   : cube_lut_3   = 14'b11101001110110;
        10'd51   : cube_lut_3   = 14'b11101001110111;
        10'd52   : cube_lut_3   = 14'b11101001111001;
        10'd53   : cube_lut_3   = 14'b11101001111010;
        10'd54   : cube_lut_3   = 14'b11101001111100;
        10'd55   : cube_lut_3   = 14'b11101001111110;
        10'd56   : cube_lut_3   = 14'b11101001111111;
        10'd57   : cube_lut_3   = 14'b11101010000001;
        10'd58   : cube_lut_3   = 14'b11101010000010;
        10'd59   : cube_lut_3   = 14'b11101010000100;
        10'd60   : cube_lut_3   = 14'b11101010000110;
        10'd61   : cube_lut_3   = 14'b11101010000111;
        10'd62   : cube_lut_3   = 14'b11101010001001;
        10'd63   : cube_lut_3   = 14'b11101010001010;
        10'd64   : cube_lut_3   = 14'b11101010001100;
        10'd65   : cube_lut_3   = 14'b11101010001110;
        10'd66   : cube_lut_3   = 14'b11101010001111;
        10'd67   : cube_lut_3   = 14'b11101010010001;
        10'd68   : cube_lut_3   = 14'b11101010010010;
        10'd69   : cube_lut_3   = 14'b11101010010100;
        10'd70   : cube_lut_3   = 14'b11101010010110;
        10'd71   : cube_lut_3   = 14'b11101010010111;
        10'd72   : cube_lut_3   = 14'b11101010011001;
        10'd73   : cube_lut_3   = 14'b11101010011010;
        10'd74   : cube_lut_3   = 14'b11101010011100;
        10'd75   : cube_lut_3   = 14'b11101010011110;
        10'd76   : cube_lut_3   = 14'b11101010011111;
        10'd77   : cube_lut_3   = 14'b11101010100001;
        10'd78   : cube_lut_3   = 14'b11101010100010;
        10'd79   : cube_lut_3   = 14'b11101010100100;
        10'd80   : cube_lut_3   = 14'b11101010100101;
        10'd81   : cube_lut_3   = 14'b11101010100111;
        10'd82   : cube_lut_3   = 14'b11101010101001;
        10'd83   : cube_lut_3   = 14'b11101010101010;
        10'd84   : cube_lut_3   = 14'b11101010101100;
        10'd85   : cube_lut_3   = 14'b11101010101101;
        10'd86   : cube_lut_3   = 14'b11101010101111;
        10'd87   : cube_lut_3   = 14'b11101010110001;
        10'd88   : cube_lut_3   = 14'b11101010110010;
        10'd89   : cube_lut_3   = 14'b11101010110100;
        10'd90   : cube_lut_3   = 14'b11101010110101;
        10'd91   : cube_lut_3   = 14'b11101010110111;
        10'd92   : cube_lut_3   = 14'b11101010111000;
        10'd93   : cube_lut_3   = 14'b11101010111010;
        10'd94   : cube_lut_3   = 14'b11101010111100;
        10'd95   : cube_lut_3   = 14'b11101010111101;
        10'd96   : cube_lut_3   = 14'b11101010111111;
        10'd97   : cube_lut_3   = 14'b11101011000000;
        10'd98   : cube_lut_3   = 14'b11101011000010;
        10'd99   : cube_lut_3   = 14'b11101011000100;
        10'd100   : cube_lut_3  = 14'b11101011000101;
        10'd101   : cube_lut_3  = 14'b11101011000111;
        10'd102   : cube_lut_3  = 14'b11101011001000;
        10'd103   : cube_lut_3  = 14'b11101011001010;
        10'd104   : cube_lut_3  = 14'b11101011001011;
        10'd105   : cube_lut_3  = 14'b11101011001101;
        10'd106   : cube_lut_3  = 14'b11101011001111;
        10'd107   : cube_lut_3  = 14'b11101011010000;
        10'd108   : cube_lut_3  = 14'b11101011010010;
        10'd109   : cube_lut_3  = 14'b11101011010011;
        10'd110   : cube_lut_3  = 14'b11101011010101;
        10'd111   : cube_lut_3  = 14'b11101011010111;
        10'd112   : cube_lut_3  = 14'b11101011011000;
        10'd113   : cube_lut_3  = 14'b11101011011010;
        10'd114   : cube_lut_3  = 14'b11101011011011;
        10'd115   : cube_lut_3  = 14'b11101011011101;
        10'd116   : cube_lut_3  = 14'b11101011011110;
        10'd117   : cube_lut_3  = 14'b11101011100000;
        10'd118   : cube_lut_3  = 14'b11101011100010;
        10'd119   : cube_lut_3  = 14'b11101011100011;
        10'd120   : cube_lut_3  = 14'b11101011100101;
        10'd121   : cube_lut_3  = 14'b11101011100110;
        10'd122   : cube_lut_3  = 14'b11101011101000;
        10'd123   : cube_lut_3  = 14'b11101011101001;
        10'd124   : cube_lut_3  = 14'b11101011101011;
        10'd125   : cube_lut_3  = 14'b11101011101101;
        10'd126   : cube_lut_3  = 14'b11101011101110;
        10'd127   : cube_lut_3  = 14'b11101011110000;
        10'd128   : cube_lut_3  = 14'b11101011110001;
        10'd129   : cube_lut_3  = 14'b11101011110011;
        10'd130   : cube_lut_3  = 14'b11101011110100;
        10'd131   : cube_lut_3  = 14'b11101011110110;
        10'd132   : cube_lut_3  = 14'b11101011111000;
        10'd133   : cube_lut_3  = 14'b11101011111001;
        10'd134   : cube_lut_3  = 14'b11101011111011;
        10'd135   : cube_lut_3  = 14'b11101011111100;
        10'd136   : cube_lut_3  = 14'b11101011111110;
        10'd137   : cube_lut_3  = 14'b11101011111111;
        10'd138   : cube_lut_3  = 14'b11101100000001;
        10'd139   : cube_lut_3  = 14'b11101100000011;
        10'd140   : cube_lut_3  = 14'b11101100000100;
        10'd141   : cube_lut_3  = 14'b11101100000110;
        10'd142   : cube_lut_3  = 14'b11101100000111;
        10'd143   : cube_lut_3  = 14'b11101100001001;
        10'd144   : cube_lut_3  = 14'b11101100001010;
        10'd145   : cube_lut_3  = 14'b11101100001100;
        10'd146   : cube_lut_3  = 14'b11101100001110;
        10'd147   : cube_lut_3  = 14'b11101100001111;
        10'd148   : cube_lut_3  = 14'b11101100010001;
        10'd149   : cube_lut_3  = 14'b11101100010010;
        10'd150   : cube_lut_3  = 14'b11101100010100;
        10'd151   : cube_lut_3  = 14'b11101100010101;
        10'd152   : cube_lut_3  = 14'b11101100010111;
        10'd153   : cube_lut_3  = 14'b11101100011000;
        10'd154   : cube_lut_3  = 14'b11101100011010;
        10'd155   : cube_lut_3  = 14'b11101100011100;
        10'd156   : cube_lut_3  = 14'b11101100011101;
        10'd157   : cube_lut_3  = 14'b11101100011111;
        10'd158   : cube_lut_3  = 14'b11101100100000;
        10'd159   : cube_lut_3  = 14'b11101100100010;
        10'd160   : cube_lut_3  = 14'b11101100100011;
        10'd161   : cube_lut_3  = 14'b11101100100101;
        10'd162   : cube_lut_3  = 14'b11101100100111;
        10'd163   : cube_lut_3  = 14'b11101100101000;
        10'd164   : cube_lut_3  = 14'b11101100101010;
        10'd165   : cube_lut_3  = 14'b11101100101011;
        10'd166   : cube_lut_3  = 14'b11101100101101;
        10'd167   : cube_lut_3  = 14'b11101100101110;
        10'd168   : cube_lut_3  = 14'b11101100110000;
        10'd169   : cube_lut_3  = 14'b11101100110001;
        10'd170   : cube_lut_3  = 14'b11101100110011;
        10'd171   : cube_lut_3  = 14'b11101100110101;
        10'd172   : cube_lut_3  = 14'b11101100110110;
        10'd173   : cube_lut_3  = 14'b11101100111000;
        10'd174   : cube_lut_3  = 14'b11101100111001;
        10'd175   : cube_lut_3  = 14'b11101100111011;
        10'd176   : cube_lut_3  = 14'b11101100111100;
        10'd177   : cube_lut_3  = 14'b11101100111110;
        10'd178   : cube_lut_3  = 14'b11101100111111;
        10'd179   : cube_lut_3  = 14'b11101101000001;
        10'd180   : cube_lut_3  = 14'b11101101000011;
        10'd181   : cube_lut_3  = 14'b11101101000100;
        10'd182   : cube_lut_3  = 14'b11101101000110;
        10'd183   : cube_lut_3  = 14'b11101101000111;
        10'd184   : cube_lut_3  = 14'b11101101001001;
        10'd185   : cube_lut_3  = 14'b11101101001010;
        10'd186   : cube_lut_3  = 14'b11101101001100;
        10'd187   : cube_lut_3  = 14'b11101101001101;
        10'd188   : cube_lut_3  = 14'b11101101001111;
        10'd189   : cube_lut_3  = 14'b11101101010001;
        10'd190   : cube_lut_3  = 14'b11101101010010;
        10'd191   : cube_lut_3  = 14'b11101101010100;
        10'd192   : cube_lut_3  = 14'b11101101010101;
        10'd193   : cube_lut_3  = 14'b11101101010111;
        10'd194   : cube_lut_3  = 14'b11101101011000;
        10'd195   : cube_lut_3  = 14'b11101101011010;
        10'd196   : cube_lut_3  = 14'b11101101011011;
        10'd197   : cube_lut_3  = 14'b11101101011101;
        10'd198   : cube_lut_3  = 14'b11101101011111;
        10'd199   : cube_lut_3  = 14'b11101101100000;
        10'd200   : cube_lut_3  = 14'b11101101100010;
        10'd201   : cube_lut_3  = 14'b11101101100011;
        10'd202   : cube_lut_3  = 14'b11101101100101;
        10'd203   : cube_lut_3  = 14'b11101101100110;
        10'd204   : cube_lut_3  = 14'b11101101101000;
        10'd205   : cube_lut_3  = 14'b11101101101001;
        10'd206   : cube_lut_3  = 14'b11101101101011;
        10'd207   : cube_lut_3  = 14'b11101101101100;
        10'd208   : cube_lut_3  = 14'b11101101101110;
        10'd209   : cube_lut_3  = 14'b11101101110000;
        10'd210   : cube_lut_3  = 14'b11101101110001;
        10'd211   : cube_lut_3  = 14'b11101101110011;
        10'd212   : cube_lut_3  = 14'b11101101110100;
        10'd213   : cube_lut_3  = 14'b11101101110110;
        10'd214   : cube_lut_3  = 14'b11101101110111;
        10'd215   : cube_lut_3  = 14'b11101101111001;
        10'd216   : cube_lut_3  = 14'b11101101111010;
        10'd217   : cube_lut_3  = 14'b11101101111100;
        10'd218   : cube_lut_3  = 14'b11101101111101;
        10'd219   : cube_lut_3  = 14'b11101101111111;
        10'd220   : cube_lut_3  = 14'b11101110000001;
        10'd221   : cube_lut_3  = 14'b11101110000010;
        10'd222   : cube_lut_3  = 14'b11101110000100;
        10'd223   : cube_lut_3  = 14'b11101110000101;
        10'd224   : cube_lut_3  = 14'b11101110000111;
        10'd225   : cube_lut_3  = 14'b11101110001000;
        10'd226   : cube_lut_3  = 14'b11101110001010;
        10'd227   : cube_lut_3  = 14'b11101110001011;
        10'd228   : cube_lut_3  = 14'b11101110001101;
        10'd229   : cube_lut_3  = 14'b11101110001110;
        10'd230   : cube_lut_3  = 14'b11101110010000;
        10'd231   : cube_lut_3  = 14'b11101110010001;
        10'd232   : cube_lut_3  = 14'b11101110010011;
        10'd233   : cube_lut_3  = 14'b11101110010101;
        10'd234   : cube_lut_3  = 14'b11101110010110;
        10'd235   : cube_lut_3  = 14'b11101110011000;
        10'd236   : cube_lut_3  = 14'b11101110011001;
        10'd237   : cube_lut_3  = 14'b11101110011011;
        10'd238   : cube_lut_3  = 14'b11101110011100;
        10'd239   : cube_lut_3  = 14'b11101110011110;
        10'd240   : cube_lut_3  = 14'b11101110011111;
        10'd241   : cube_lut_3  = 14'b11101110100001;
        10'd242   : cube_lut_3  = 14'b11101110100010;
        10'd243   : cube_lut_3  = 14'b11101110100100;
        10'd244   : cube_lut_3  = 14'b11101110100101;
        10'd245   : cube_lut_3  = 14'b11101110100111;
        10'd246   : cube_lut_3  = 14'b11101110101001;
        10'd247   : cube_lut_3  = 14'b11101110101010;
        10'd248   : cube_lut_3  = 14'b11101110101100;
        10'd249   : cube_lut_3  = 14'b11101110101101;
        10'd250   : cube_lut_3  = 14'b11101110101111;
        10'd251   : cube_lut_3  = 14'b11101110110000;
        10'd252   : cube_lut_3  = 14'b11101110110010;
        10'd253   : cube_lut_3  = 14'b11101110110011;
        10'd254   : cube_lut_3  = 14'b11101110110101;
        10'd255   : cube_lut_3  = 14'b11101110110110;
        10'd256   : cube_lut_3  = 14'b11101110111000;
        10'd257   : cube_lut_3  = 14'b11101110111001;
        10'd258   : cube_lut_3  = 14'b11101110111011;
        10'd259   : cube_lut_3  = 14'b11101110111100;
        10'd260   : cube_lut_3  = 14'b11101110111110;
        10'd261   : cube_lut_3  = 14'b11101111000000;
        10'd262   : cube_lut_3  = 14'b11101111000001;
        10'd263   : cube_lut_3  = 14'b11101111000011;
        10'd264   : cube_lut_3  = 14'b11101111000100;
        10'd265   : cube_lut_3  = 14'b11101111000110;
        10'd266   : cube_lut_3  = 14'b11101111000111;
        10'd267   : cube_lut_3  = 14'b11101111001001;
        10'd268   : cube_lut_3  = 14'b11101111001010;
        10'd269   : cube_lut_3  = 14'b11101111001100;
        10'd270   : cube_lut_3  = 14'b11101111001101;
        10'd271   : cube_lut_3  = 14'b11101111001111;
        10'd272   : cube_lut_3  = 14'b11101111010000;
        10'd273   : cube_lut_3  = 14'b11101111010010;
        10'd274   : cube_lut_3  = 14'b11101111010011;
        10'd275   : cube_lut_3  = 14'b11101111010101;
        10'd276   : cube_lut_3  = 14'b11101111010110;
        10'd277   : cube_lut_3  = 14'b11101111011000;
        10'd278   : cube_lut_3  = 14'b11101111011001;
        10'd279   : cube_lut_3  = 14'b11101111011011;
        10'd280   : cube_lut_3  = 14'b11101111011101;
        10'd281   : cube_lut_3  = 14'b11101111011110;
        10'd282   : cube_lut_3  = 14'b11101111100000;
        10'd283   : cube_lut_3  = 14'b11101111100001;
        10'd284   : cube_lut_3  = 14'b11101111100011;
        10'd285   : cube_lut_3  = 14'b11101111100100;
        10'd286   : cube_lut_3  = 14'b11101111100110;
        10'd287   : cube_lut_3  = 14'b11101111100111;
        10'd288   : cube_lut_3  = 14'b11101111101001;
        10'd289   : cube_lut_3  = 14'b11101111101010;
        10'd290   : cube_lut_3  = 14'b11101111101100;
        10'd291   : cube_lut_3  = 14'b11101111101101;
        10'd292   : cube_lut_3  = 14'b11101111101111;
        10'd293   : cube_lut_3  = 14'b11101111110000;
        10'd294   : cube_lut_3  = 14'b11101111110010;
        10'd295   : cube_lut_3  = 14'b11101111110011;
        10'd296   : cube_lut_3  = 14'b11101111110101;
        10'd297   : cube_lut_3  = 14'b11101111110110;
        10'd298   : cube_lut_3  = 14'b11101111111000;
        10'd299   : cube_lut_3  = 14'b11101111111001;
        10'd300   : cube_lut_3  = 14'b11101111111011;
        10'd301   : cube_lut_3  = 14'b11101111111100;
        10'd302   : cube_lut_3  = 14'b11101111111110;
        10'd303   : cube_lut_3  = 14'b11110000000000;
        10'd304   : cube_lut_3  = 14'b11110000000001;
        10'd305   : cube_lut_3  = 14'b11110000000011;
        10'd306   : cube_lut_3  = 14'b11110000000100;
        10'd307   : cube_lut_3  = 14'b11110000000110;
        10'd308   : cube_lut_3  = 14'b11110000000111;
        10'd309   : cube_lut_3  = 14'b11110000001001;
        10'd310   : cube_lut_3  = 14'b11110000001010;
        10'd311   : cube_lut_3  = 14'b11110000001100;
        10'd312   : cube_lut_3  = 14'b11110000001101;
        10'd313   : cube_lut_3  = 14'b11110000001111;
        10'd314   : cube_lut_3  = 14'b11110000010000;
        10'd315   : cube_lut_3  = 14'b11110000010010;
        10'd316   : cube_lut_3  = 14'b11110000010011;
        10'd317   : cube_lut_3  = 14'b11110000010101;
        10'd318   : cube_lut_3  = 14'b11110000010110;
        10'd319   : cube_lut_3  = 14'b11110000011000;
        10'd320   : cube_lut_3  = 14'b11110000011001;
        10'd321   : cube_lut_3  = 14'b11110000011011;
        10'd322   : cube_lut_3  = 14'b11110000011100;
        10'd323   : cube_lut_3  = 14'b11110000011110;
        10'd324   : cube_lut_3  = 14'b11110000011111;
        10'd325   : cube_lut_3  = 14'b11110000100001;
        10'd326   : cube_lut_3  = 14'b11110000100010;
        10'd327   : cube_lut_3  = 14'b11110000100100;
        10'd328   : cube_lut_3  = 14'b11110000100101;
        10'd329   : cube_lut_3  = 14'b11110000100111;
        10'd330   : cube_lut_3  = 14'b11110000101000;
        10'd331   : cube_lut_3  = 14'b11110000101010;
        10'd332   : cube_lut_3  = 14'b11110000101011;
        10'd333   : cube_lut_3  = 14'b11110000101101;
        10'd334   : cube_lut_3  = 14'b11110000101110;
        10'd335   : cube_lut_3  = 14'b11110000110000;
        10'd336   : cube_lut_3  = 14'b11110000110001;
        10'd337   : cube_lut_3  = 14'b11110000110011;
        10'd338   : cube_lut_3  = 14'b11110000110100;
        10'd339   : cube_lut_3  = 14'b11110000110110;
        10'd340   : cube_lut_3  = 14'b11110000110111;
        10'd341   : cube_lut_3  = 14'b11110000111001;
        10'd342   : cube_lut_3  = 14'b11110000111010;
        10'd343   : cube_lut_3  = 14'b11110000111100;
        10'd344   : cube_lut_3  = 14'b11110000111101;
        10'd345   : cube_lut_3  = 14'b11110000111111;
        10'd346   : cube_lut_3  = 14'b11110001000000;
        10'd347   : cube_lut_3  = 14'b11110001000010;
        10'd348   : cube_lut_3  = 14'b11110001000011;
        10'd349   : cube_lut_3  = 14'b11110001000101;
        10'd350   : cube_lut_3  = 14'b11110001000110;
        10'd351   : cube_lut_3  = 14'b11110001001000;
        10'd352   : cube_lut_3  = 14'b11110001001001;
        10'd353   : cube_lut_3  = 14'b11110001001011;
        10'd354   : cube_lut_3  = 14'b11110001001100;
        10'd355   : cube_lut_3  = 14'b11110001001110;
        10'd356   : cube_lut_3  = 14'b11110001001111;
        10'd357   : cube_lut_3  = 14'b11110001010001;
        10'd358   : cube_lut_3  = 14'b11110001010010;
        10'd359   : cube_lut_3  = 14'b11110001010100;
        10'd360   : cube_lut_3  = 14'b11110001010101;
        10'd361   : cube_lut_3  = 14'b11110001010111;
        10'd362   : cube_lut_3  = 14'b11110001011000;
        10'd363   : cube_lut_3  = 14'b11110001011010;
        10'd364   : cube_lut_3  = 14'b11110001011011;
        10'd365   : cube_lut_3  = 14'b11110001011101;
        10'd366   : cube_lut_3  = 14'b11110001011110;
        10'd367   : cube_lut_3  = 14'b11110001100000;
        10'd368   : cube_lut_3  = 14'b11110001100001;
        10'd369   : cube_lut_3  = 14'b11110001100011;
        10'd370   : cube_lut_3  = 14'b11110001100100;
        10'd371   : cube_lut_3  = 14'b11110001100110;
        10'd372   : cube_lut_3  = 14'b11110001100111;
        10'd373   : cube_lut_3  = 14'b11110001101001;
        10'd374   : cube_lut_3  = 14'b11110001101010;
        10'd375   : cube_lut_3  = 14'b11110001101100;
        10'd376   : cube_lut_3  = 14'b11110001101101;
        10'd377   : cube_lut_3  = 14'b11110001101111;
        10'd378   : cube_lut_3  = 14'b11110001110000;
        10'd379   : cube_lut_3  = 14'b11110001110010;
        10'd380   : cube_lut_3  = 14'b11110001110011;
        10'd381   : cube_lut_3  = 14'b11110001110101;
        10'd382   : cube_lut_3  = 14'b11110001110110;
        10'd383   : cube_lut_3  = 14'b11110001111000;
        10'd384   : cube_lut_3  = 14'b11110001111001;
        10'd385   : cube_lut_3  = 14'b11110001111011;
        10'd386   : cube_lut_3  = 14'b11110001111100;
        10'd387   : cube_lut_3  = 14'b11110001111110;
        10'd388   : cube_lut_3  = 14'b11110001111111;
        10'd389   : cube_lut_3  = 14'b11110010000001;
        10'd390   : cube_lut_3  = 14'b11110010000010;
        10'd391   : cube_lut_3  = 14'b11110010000100;
        10'd392   : cube_lut_3  = 14'b11110010000101;
        10'd393   : cube_lut_3  = 14'b11110010000111;
        10'd394   : cube_lut_3  = 14'b11110010001000;
        10'd395   : cube_lut_3  = 14'b11110010001010;
        10'd396   : cube_lut_3  = 14'b11110010001011;
        10'd397   : cube_lut_3  = 14'b11110010001101;
        10'd398   : cube_lut_3  = 14'b11110010001110;
        10'd399   : cube_lut_3  = 14'b11110010010000;
        10'd400   : cube_lut_3  = 14'b11110010010001;
        10'd401   : cube_lut_3  = 14'b11110010010011;
        10'd402   : cube_lut_3  = 14'b11110010010100;
        10'd403   : cube_lut_3  = 14'b11110010010110;
        10'd404   : cube_lut_3  = 14'b11110010010111;
        10'd405   : cube_lut_3  = 14'b11110010011001;
        10'd406   : cube_lut_3  = 14'b11110010011010;
        10'd407   : cube_lut_3  = 14'b11110010011100;
        10'd408   : cube_lut_3  = 14'b11110010011101;
        10'd409   : cube_lut_3  = 14'b11110010011111;
        10'd410   : cube_lut_3  = 14'b11110010100000;
        10'd411   : cube_lut_3  = 14'b11110010100010;
        10'd412   : cube_lut_3  = 14'b11110010100011;
        10'd413   : cube_lut_3  = 14'b11110010100101;
        10'd414   : cube_lut_3  = 14'b11110010100110;
        10'd415   : cube_lut_3  = 14'b11110010101000;
        10'd416   : cube_lut_3  = 14'b11110010101001;
        10'd417   : cube_lut_3  = 14'b11110010101011;
        10'd418   : cube_lut_3  = 14'b11110010101100;
        10'd419   : cube_lut_3  = 14'b11110010101101;
        10'd420   : cube_lut_3  = 14'b11110010101111;
        10'd421   : cube_lut_3  = 14'b11110010110000;
        10'd422   : cube_lut_3  = 14'b11110010110010;
        10'd423   : cube_lut_3  = 14'b11110010110011;
        10'd424   : cube_lut_3  = 14'b11110010110101;
        10'd425   : cube_lut_3  = 14'b11110010110110;
        10'd426   : cube_lut_3  = 14'b11110010111000;
        10'd427   : cube_lut_3  = 14'b11110010111001;
        10'd428   : cube_lut_3  = 14'b11110010111011;
        10'd429   : cube_lut_3  = 14'b11110010111100;
        10'd430   : cube_lut_3  = 14'b11110010111110;
        10'd431   : cube_lut_3  = 14'b11110010111111;
        10'd432   : cube_lut_3  = 14'b11110011000001;
        10'd433   : cube_lut_3  = 14'b11110011000010;
        10'd434   : cube_lut_3  = 14'b11110011000100;
        10'd435   : cube_lut_3  = 14'b11110011000101;
        10'd436   : cube_lut_3  = 14'b11110011000111;
        10'd437   : cube_lut_3  = 14'b11110011001000;
        10'd438   : cube_lut_3  = 14'b11110011001010;
        10'd439   : cube_lut_3  = 14'b11110011001011;
        10'd440   : cube_lut_3  = 14'b11110011001101;
        10'd441   : cube_lut_3  = 14'b11110011001110;
        10'd442   : cube_lut_3  = 14'b11110011010000;
        10'd443   : cube_lut_3  = 14'b11110011010001;
        10'd444   : cube_lut_3  = 14'b11110011010010;
        10'd445   : cube_lut_3  = 14'b11110011010100;
        10'd446   : cube_lut_3  = 14'b11110011010101;
        10'd447   : cube_lut_3  = 14'b11110011010111;
        10'd448   : cube_lut_3  = 14'b11110011011000;
        10'd449   : cube_lut_3  = 14'b11110011011010;
        10'd450   : cube_lut_3  = 14'b11110011011011;
        10'd451   : cube_lut_3  = 14'b11110011011101;
        10'd452   : cube_lut_3  = 14'b11110011011110;
        10'd453   : cube_lut_3  = 14'b11110011100000;
        10'd454   : cube_lut_3  = 14'b11110011100001;
        10'd455   : cube_lut_3  = 14'b11110011100011;
        10'd456   : cube_lut_3  = 14'b11110011100100;
        10'd457   : cube_lut_3  = 14'b11110011100110;
        10'd458   : cube_lut_3  = 14'b11110011100111;
        10'd459   : cube_lut_3  = 14'b11110011101001;
        10'd460   : cube_lut_3  = 14'b11110011101010;
        10'd461   : cube_lut_3  = 14'b11110011101100;
        10'd462   : cube_lut_3  = 14'b11110011101101;
        10'd463   : cube_lut_3  = 14'b11110011101110;
        10'd464   : cube_lut_3  = 14'b11110011110000;
        10'd465   : cube_lut_3  = 14'b11110011110001;
        10'd466   : cube_lut_3  = 14'b11110011110011;
        10'd467   : cube_lut_3  = 14'b11110011110100;
        10'd468   : cube_lut_3  = 14'b11110011110110;
        10'd469   : cube_lut_3  = 14'b11110011110111;
        10'd470   : cube_lut_3  = 14'b11110011111001;
        10'd471   : cube_lut_3  = 14'b11110011111010;
        10'd472   : cube_lut_3  = 14'b11110011111100;
        10'd473   : cube_lut_3  = 14'b11110011111101;
        10'd474   : cube_lut_3  = 14'b11110011111111;
        10'd475   : cube_lut_3  = 14'b11110100000000;
        10'd476   : cube_lut_3  = 14'b11110100000010;
        10'd477   : cube_lut_3  = 14'b11110100000011;
        10'd478   : cube_lut_3  = 14'b11110100000101;
        10'd479   : cube_lut_3  = 14'b11110100000110;
        10'd480   : cube_lut_3  = 14'b11110100000111;
        10'd481   : cube_lut_3  = 14'b11110100001001;
        10'd482   : cube_lut_3  = 14'b11110100001010;
        10'd483   : cube_lut_3  = 14'b11110100001100;
        10'd484   : cube_lut_3  = 14'b11110100001101;
        10'd485   : cube_lut_3  = 14'b11110100001111;
        10'd486   : cube_lut_3  = 14'b11110100010000;
        10'd487   : cube_lut_3  = 14'b11110100010010;
        10'd488   : cube_lut_3  = 14'b11110100010011;
        10'd489   : cube_lut_3  = 14'b11110100010101;
        10'd490   : cube_lut_3  = 14'b11110100010110;
        10'd491   : cube_lut_3  = 14'b11110100011000;
        10'd492   : cube_lut_3  = 14'b11110100011001;
        10'd493   : cube_lut_3  = 14'b11110100011010;
        10'd494   : cube_lut_3  = 14'b11110100011100;
        10'd495   : cube_lut_3  = 14'b11110100011101;
        10'd496   : cube_lut_3  = 14'b11110100011111;
        10'd497   : cube_lut_3  = 14'b11110100100000;
        10'd498   : cube_lut_3  = 14'b11110100100010;
        10'd499   : cube_lut_3  = 14'b11110100100011;
        10'd500   : cube_lut_3  = 14'b11110100100101;
        10'd501   : cube_lut_3  = 14'b11110100100110;
        10'd502   : cube_lut_3  = 14'b11110100101000;
        10'd503   : cube_lut_3  = 14'b11110100101001;
        10'd504   : cube_lut_3  = 14'b11110100101011;
        10'd505   : cube_lut_3  = 14'b11110100101100;
        10'd506   : cube_lut_3  = 14'b11110100101101;
        10'd507   : cube_lut_3  = 14'b11110100101111;
        10'd508   : cube_lut_3  = 14'b11110100110000;
        10'd509   : cube_lut_3  = 14'b11110100110010;
        10'd510   : cube_lut_3  = 14'b11110100110011;
        10'd511   : cube_lut_3  = 14'b11110100110101;
        10'd512   : cube_lut_3  = 14'b11110100110110;
        10'd513   : cube_lut_3  = 14'b11110100111000;
        10'd514   : cube_lut_3  = 14'b11110100111001;
        10'd515   : cube_lut_3  = 14'b11110100111011;
        10'd516   : cube_lut_3  = 14'b11110100111100;
        10'd517   : cube_lut_3  = 14'b11110100111110;
        10'd518   : cube_lut_3  = 14'b11110100111111;
        10'd519   : cube_lut_3  = 14'b11110101000000;
        10'd520   : cube_lut_3  = 14'b11110101000010;
        10'd521   : cube_lut_3  = 14'b11110101000011;
        10'd522   : cube_lut_3  = 14'b11110101000101;
        10'd523   : cube_lut_3  = 14'b11110101000110;
        10'd524   : cube_lut_3  = 14'b11110101001000;
        10'd525   : cube_lut_3  = 14'b11110101001001;
        10'd526   : cube_lut_3  = 14'b11110101001011;
        10'd527   : cube_lut_3  = 14'b11110101001100;
        10'd528   : cube_lut_3  = 14'b11110101001110;
        10'd529   : cube_lut_3  = 14'b11110101001111;
        10'd530   : cube_lut_3  = 14'b11110101010000;
        10'd531   : cube_lut_3  = 14'b11110101010010;
        10'd532   : cube_lut_3  = 14'b11110101010011;
        10'd533   : cube_lut_3  = 14'b11110101010101;
        10'd534   : cube_lut_3  = 14'b11110101010110;
        10'd535   : cube_lut_3  = 14'b11110101011000;
        10'd536   : cube_lut_3  = 14'b11110101011001;
        10'd537   : cube_lut_3  = 14'b11110101011011;
        10'd538   : cube_lut_3  = 14'b11110101011100;
        10'd539   : cube_lut_3  = 14'b11110101011101;
        10'd540   : cube_lut_3  = 14'b11110101011111;
        10'd541   : cube_lut_3  = 14'b11110101100000;
        10'd542   : cube_lut_3  = 14'b11110101100010;
        10'd543   : cube_lut_3  = 14'b11110101100011;
        10'd544   : cube_lut_3  = 14'b11110101100101;
        10'd545   : cube_lut_3  = 14'b11110101100110;
        10'd546   : cube_lut_3  = 14'b11110101101000;
        10'd547   : cube_lut_3  = 14'b11110101101001;
        10'd548   : cube_lut_3  = 14'b11110101101011;
        10'd549   : cube_lut_3  = 14'b11110101101100;
        10'd550   : cube_lut_3  = 14'b11110101101101;
        10'd551   : cube_lut_3  = 14'b11110101101111;
        10'd552   : cube_lut_3  = 14'b11110101110000;
        10'd553   : cube_lut_3  = 14'b11110101110010;
        10'd554   : cube_lut_3  = 14'b11110101110011;
        10'd555   : cube_lut_3  = 14'b11110101110101;
        10'd556   : cube_lut_3  = 14'b11110101110110;
        10'd557   : cube_lut_3  = 14'b11110101111000;
        10'd558   : cube_lut_3  = 14'b11110101111001;
        10'd559   : cube_lut_3  = 14'b11110101111010;
        10'd560   : cube_lut_3  = 14'b11110101111100;
        10'd561   : cube_lut_3  = 14'b11110101111101;
        10'd562   : cube_lut_3  = 14'b11110101111111;
        10'd563   : cube_lut_3  = 14'b11110110000000;
        10'd564   : cube_lut_3  = 14'b11110110000010;
        10'd565   : cube_lut_3  = 14'b11110110000011;
        10'd566   : cube_lut_3  = 14'b11110110000101;
        10'd567   : cube_lut_3  = 14'b11110110000110;
        10'd568   : cube_lut_3  = 14'b11110110000111;
        10'd569   : cube_lut_3  = 14'b11110110001001;
        10'd570   : cube_lut_3  = 14'b11110110001010;
        10'd571   : cube_lut_3  = 14'b11110110001100;
        10'd572   : cube_lut_3  = 14'b11110110001101;
        10'd573   : cube_lut_3  = 14'b11110110001111;
        10'd574   : cube_lut_3  = 14'b11110110010000;
        10'd575   : cube_lut_3  = 14'b11110110010010;
        10'd576   : cube_lut_3  = 14'b11110110010011;
        10'd577   : cube_lut_3  = 14'b11110110010100;
        10'd578   : cube_lut_3  = 14'b11110110010110;
        10'd579   : cube_lut_3  = 14'b11110110010111;
        10'd580   : cube_lut_3  = 14'b11110110011001;
        10'd581   : cube_lut_3  = 14'b11110110011010;
        10'd582   : cube_lut_3  = 14'b11110110011100;
        10'd583   : cube_lut_3  = 14'b11110110011101;
        10'd584   : cube_lut_3  = 14'b11110110011110;
        10'd585   : cube_lut_3  = 14'b11110110100000;
        10'd586   : cube_lut_3  = 14'b11110110100001;
        10'd587   : cube_lut_3  = 14'b11110110100011;
        10'd588   : cube_lut_3  = 14'b11110110100100;
        10'd589   : cube_lut_3  = 14'b11110110100110;
        10'd590   : cube_lut_3  = 14'b11110110100111;
        10'd591   : cube_lut_3  = 14'b11110110101001;
        10'd592   : cube_lut_3  = 14'b11110110101010;
        10'd593   : cube_lut_3  = 14'b11110110101011;
        10'd594   : cube_lut_3  = 14'b11110110101101;
        10'd595   : cube_lut_3  = 14'b11110110101110;
        10'd596   : cube_lut_3  = 14'b11110110110000;
        10'd597   : cube_lut_3  = 14'b11110110110001;
        10'd598   : cube_lut_3  = 14'b11110110110011;
        10'd599   : cube_lut_3  = 14'b11110110110100;
        10'd600   : cube_lut_3  = 14'b11110110110101;
        10'd601   : cube_lut_3  = 14'b11110110110111;
        10'd602   : cube_lut_3  = 14'b11110110111000;
        10'd603   : cube_lut_3  = 14'b11110110111010;
        10'd604   : cube_lut_3  = 14'b11110110111011;
        10'd605   : cube_lut_3  = 14'b11110110111101;
        10'd606   : cube_lut_3  = 14'b11110110111110;
        10'd607   : cube_lut_3  = 14'b11110110111111;
        10'd608   : cube_lut_3  = 14'b11110111000001;
        10'd609   : cube_lut_3  = 14'b11110111000010;
        10'd610   : cube_lut_3  = 14'b11110111000100;
        10'd611   : cube_lut_3  = 14'b11110111000101;
        10'd612   : cube_lut_3  = 14'b11110111000111;
        10'd613   : cube_lut_3  = 14'b11110111001000;
        10'd614   : cube_lut_3  = 14'b11110111001010;
        10'd615   : cube_lut_3  = 14'b11110111001011;
        10'd616   : cube_lut_3  = 14'b11110111001100;
        10'd617   : cube_lut_3  = 14'b11110111001110;
        10'd618   : cube_lut_3  = 14'b11110111001111;
        10'd619   : cube_lut_3  = 14'b11110111010001;
        10'd620   : cube_lut_3  = 14'b11110111010010;
        10'd621   : cube_lut_3  = 14'b11110111010100;
        10'd622   : cube_lut_3  = 14'b11110111010101;
        10'd623   : cube_lut_3  = 14'b11110111010110;
        10'd624   : cube_lut_3  = 14'b11110111011000;
        10'd625   : cube_lut_3  = 14'b11110111011001;
        10'd626   : cube_lut_3  = 14'b11110111011011;
        10'd627   : cube_lut_3  = 14'b11110111011100;
        10'd628   : cube_lut_3  = 14'b11110111011110;
        10'd629   : cube_lut_3  = 14'b11110111011111;
        10'd630   : cube_lut_3  = 14'b11110111100000;
        10'd631   : cube_lut_3  = 14'b11110111100010;
        10'd632   : cube_lut_3  = 14'b11110111100011;
        10'd633   : cube_lut_3  = 14'b11110111100101;
        10'd634   : cube_lut_3  = 14'b11110111100110;
        10'd635   : cube_lut_3  = 14'b11110111100111;
        10'd636   : cube_lut_3  = 14'b11110111101001;
        10'd637   : cube_lut_3  = 14'b11110111101010;
        10'd638   : cube_lut_3  = 14'b11110111101100;
        10'd639   : cube_lut_3  = 14'b11110111101101;
        10'd640   : cube_lut_3  = 14'b11110111101111;
        10'd641   : cube_lut_3  = 14'b11110111110000;
        10'd642   : cube_lut_3  = 14'b11110111110001;
        10'd643   : cube_lut_3  = 14'b11110111110011;
        10'd644   : cube_lut_3  = 14'b11110111110100;
        10'd645   : cube_lut_3  = 14'b11110111110110;
        10'd646   : cube_lut_3  = 14'b11110111110111;
        10'd647   : cube_lut_3  = 14'b11110111111001;
        10'd648   : cube_lut_3  = 14'b11110111111010;
        10'd649   : cube_lut_3  = 14'b11110111111011;
        10'd650   : cube_lut_3  = 14'b11110111111101;
        10'd651   : cube_lut_3  = 14'b11110111111110;
        10'd652   : cube_lut_3  = 14'b11111000000000;
        10'd653   : cube_lut_3  = 14'b11111000000001;
        10'd654   : cube_lut_3  = 14'b11111000000011;
        10'd655   : cube_lut_3  = 14'b11111000000100;
        10'd656   : cube_lut_3  = 14'b11111000000101;
        10'd657   : cube_lut_3  = 14'b11111000000111;
        10'd658   : cube_lut_3  = 14'b11111000001000;
        10'd659   : cube_lut_3  = 14'b11111000001010;
        10'd660   : cube_lut_3  = 14'b11111000001011;
        10'd661   : cube_lut_3  = 14'b11111000001100;
        10'd662   : cube_lut_3  = 14'b11111000001110;
        10'd663   : cube_lut_3  = 14'b11111000001111;
        10'd664   : cube_lut_3  = 14'b11111000010001;
        10'd665   : cube_lut_3  = 14'b11111000010010;
        10'd666   : cube_lut_3  = 14'b11111000010100;
        10'd667   : cube_lut_3  = 14'b11111000010101;
        10'd668   : cube_lut_3  = 14'b11111000010110;
        10'd669   : cube_lut_3  = 14'b11111000011000;
        10'd670   : cube_lut_3  = 14'b11111000011001;
        10'd671   : cube_lut_3  = 14'b11111000011011;
        10'd672   : cube_lut_3  = 14'b11111000011100;
        10'd673   : cube_lut_3  = 14'b11111000011101;
        10'd674   : cube_lut_3  = 14'b11111000011111;
        10'd675   : cube_lut_3  = 14'b11111000100000;
        10'd676   : cube_lut_3  = 14'b11111000100010;
        10'd677   : cube_lut_3  = 14'b11111000100011;
        10'd678   : cube_lut_3  = 14'b11111000100101;
        10'd679   : cube_lut_3  = 14'b11111000100110;
        10'd680   : cube_lut_3  = 14'b11111000100111;
        10'd681   : cube_lut_3  = 14'b11111000101001;
        10'd682   : cube_lut_3  = 14'b11111000101010;
        10'd683   : cube_lut_3  = 14'b11111000101100;
        10'd684   : cube_lut_3  = 14'b11111000101101;
        10'd685   : cube_lut_3  = 14'b11111000101110;
        10'd686   : cube_lut_3  = 14'b11111000110000;
        10'd687   : cube_lut_3  = 14'b11111000110001;
        10'd688   : cube_lut_3  = 14'b11111000110011;
        10'd689   : cube_lut_3  = 14'b11111000110100;
        10'd690   : cube_lut_3  = 14'b11111000110101;
        10'd691   : cube_lut_3  = 14'b11111000110111;
        10'd692   : cube_lut_3  = 14'b11111000111000;
        10'd693   : cube_lut_3  = 14'b11111000111010;
        10'd694   : cube_lut_3  = 14'b11111000111011;
        10'd695   : cube_lut_3  = 14'b11111000111101;
        10'd696   : cube_lut_3  = 14'b11111000111110;
        10'd697   : cube_lut_3  = 14'b11111000111111;
        10'd698   : cube_lut_3  = 14'b11111001000001;
        10'd699   : cube_lut_3  = 14'b11111001000010;
        10'd700   : cube_lut_3  = 14'b11111001000100;
        10'd701   : cube_lut_3  = 14'b11111001000101;
        10'd702   : cube_lut_3  = 14'b11111001000110;
        10'd703   : cube_lut_3  = 14'b11111001001000;
        10'd704   : cube_lut_3  = 14'b11111001001001;
        10'd705   : cube_lut_3  = 14'b11111001001011;
        10'd706   : cube_lut_3  = 14'b11111001001100;
        10'd707   : cube_lut_3  = 14'b11111001001101;
        10'd708   : cube_lut_3  = 14'b11111001001111;
        10'd709   : cube_lut_3  = 14'b11111001010000;
        10'd710   : cube_lut_3  = 14'b11111001010010;
        10'd711   : cube_lut_3  = 14'b11111001010011;
        10'd712   : cube_lut_3  = 14'b11111001010100;
        10'd713   : cube_lut_3  = 14'b11111001010110;
        10'd714   : cube_lut_3  = 14'b11111001010111;
        10'd715   : cube_lut_3  = 14'b11111001011001;
        10'd716   : cube_lut_3  = 14'b11111001011010;
        10'd717   : cube_lut_3  = 14'b11111001011011;
        10'd718   : cube_lut_3  = 14'b11111001011101;
        10'd719   : cube_lut_3  = 14'b11111001011110;
        10'd720   : cube_lut_3  = 14'b11111001100000;
        10'd721   : cube_lut_3  = 14'b11111001100001;
        10'd722   : cube_lut_3  = 14'b11111001100011;
        10'd723   : cube_lut_3  = 14'b11111001100100;
        10'd724   : cube_lut_3  = 14'b11111001100101;
        10'd725   : cube_lut_3  = 14'b11111001100111;
        10'd726   : cube_lut_3  = 14'b11111001101000;
        10'd727   : cube_lut_3  = 14'b11111001101010;
        10'd728   : cube_lut_3  = 14'b11111001101011;
        10'd729   : cube_lut_3  = 14'b11111001101100;
        10'd730   : cube_lut_3  = 14'b11111001101110;
        10'd731   : cube_lut_3  = 14'b11111001101111;
        10'd732   : cube_lut_3  = 14'b11111001110001;
        10'd733   : cube_lut_3  = 14'b11111001110010;
        10'd734   : cube_lut_3  = 14'b11111001110011;
        10'd735   : cube_lut_3  = 14'b11111001110101;
        10'd736   : cube_lut_3  = 14'b11111001110110;
        10'd737   : cube_lut_3  = 14'b11111001111000;
        10'd738   : cube_lut_3  = 14'b11111001111001;
        10'd739   : cube_lut_3  = 14'b11111001111010;
        10'd740   : cube_lut_3  = 14'b11111001111100;
        10'd741   : cube_lut_3  = 14'b11111001111101;
        10'd742   : cube_lut_3  = 14'b11111001111111;
        10'd743   : cube_lut_3  = 14'b11111010000000;
        10'd744   : cube_lut_3  = 14'b11111010000001;
        10'd745   : cube_lut_3  = 14'b11111010000011;
        10'd746   : cube_lut_3  = 14'b11111010000100;
        10'd747   : cube_lut_3  = 14'b11111010000110;
        10'd748   : cube_lut_3  = 14'b11111010000111;
        10'd749   : cube_lut_3  = 14'b11111010001000;
        10'd750   : cube_lut_3  = 14'b11111010001010;
        10'd751   : cube_lut_3  = 14'b11111010001011;
        10'd752   : cube_lut_3  = 14'b11111010001100;
        10'd753   : cube_lut_3  = 14'b11111010001110;
        10'd754   : cube_lut_3  = 14'b11111010001111;
        10'd755   : cube_lut_3  = 14'b11111010010001;
        10'd756   : cube_lut_3  = 14'b11111010010010;
        10'd757   : cube_lut_3  = 14'b11111010010011;
        10'd758   : cube_lut_3  = 14'b11111010010101;
        10'd759   : cube_lut_3  = 14'b11111010010110;
        10'd760   : cube_lut_3  = 14'b11111010011000;
        10'd761   : cube_lut_3  = 14'b11111010011001;
        10'd762   : cube_lut_3  = 14'b11111010011010;
        10'd763   : cube_lut_3  = 14'b11111010011100;
        10'd764   : cube_lut_3  = 14'b11111010011101;
        10'd765   : cube_lut_3  = 14'b11111010011111;
        10'd766   : cube_lut_3  = 14'b11111010100000;
        10'd767   : cube_lut_3  = 14'b11111010100001;
        10'd768   : cube_lut_3  = 14'b11111010100011;
        10'd769   : cube_lut_3  = 14'b11111010100100;
        10'd770   : cube_lut_3  = 14'b11111010100110;
        10'd771   : cube_lut_3  = 14'b11111010100111;
        10'd772   : cube_lut_3  = 14'b11111010101000;
        10'd773   : cube_lut_3  = 14'b11111010101010;
        10'd774   : cube_lut_3  = 14'b11111010101011;
        10'd775   : cube_lut_3  = 14'b11111010101101;
        10'd776   : cube_lut_3  = 14'b11111010101110;
        10'd777   : cube_lut_3  = 14'b11111010101111;
        10'd778   : cube_lut_3  = 14'b11111010110001;
        10'd779   : cube_lut_3  = 14'b11111010110010;
        10'd780   : cube_lut_3  = 14'b11111010110011;
        10'd781   : cube_lut_3  = 14'b11111010110101;
        10'd782   : cube_lut_3  = 14'b11111010110110;
        10'd783   : cube_lut_3  = 14'b11111010111000;
        10'd784   : cube_lut_3  = 14'b11111010111001;
        10'd785   : cube_lut_3  = 14'b11111010111010;
        10'd786   : cube_lut_3  = 14'b11111010111100;
        10'd787   : cube_lut_3  = 14'b11111010111101;
        10'd788   : cube_lut_3  = 14'b11111010111111;
        10'd789   : cube_lut_3  = 14'b11111011000000;
        10'd790   : cube_lut_3  = 14'b11111011000001;
        10'd791   : cube_lut_3  = 14'b11111011000011;
        10'd792   : cube_lut_3  = 14'b11111011000100;
        10'd793   : cube_lut_3  = 14'b11111011000110;
        10'd794   : cube_lut_3  = 14'b11111011000111;
        10'd795   : cube_lut_3  = 14'b11111011001000;
        10'd796   : cube_lut_3  = 14'b11111011001010;
        10'd797   : cube_lut_3  = 14'b11111011001011;
        10'd798   : cube_lut_3  = 14'b11111011001100;
        10'd799   : cube_lut_3  = 14'b11111011001110;
        10'd800   : cube_lut_3  = 14'b11111011001111;
        10'd801   : cube_lut_3  = 14'b11111011010001;
        10'd802   : cube_lut_3  = 14'b11111011010010;
        10'd803   : cube_lut_3  = 14'b11111011010011;
        10'd804   : cube_lut_3  = 14'b11111011010101;
        10'd805   : cube_lut_3  = 14'b11111011010110;
        10'd806   : cube_lut_3  = 14'b11111011011000;
        10'd807   : cube_lut_3  = 14'b11111011011001;
        10'd808   : cube_lut_3  = 14'b11111011011010;
        10'd809   : cube_lut_3  = 14'b11111011011100;
        10'd810   : cube_lut_3  = 14'b11111011011101;
        10'd811   : cube_lut_3  = 14'b11111011011110;
        10'd812   : cube_lut_3  = 14'b11111011100000;
        10'd813   : cube_lut_3  = 14'b11111011100001;
        10'd814   : cube_lut_3  = 14'b11111011100011;
        10'd815   : cube_lut_3  = 14'b11111011100100;
        10'd816   : cube_lut_3  = 14'b11111011100101;
        10'd817   : cube_lut_3  = 14'b11111011100111;
        10'd818   : cube_lut_3  = 14'b11111011101000;
        10'd819   : cube_lut_3  = 14'b11111011101001;
        10'd820   : cube_lut_3  = 14'b11111011101011;
        10'd821   : cube_lut_3  = 14'b11111011101100;
        10'd822   : cube_lut_3  = 14'b11111011101110;
        10'd823   : cube_lut_3  = 14'b11111011101111;
        10'd824   : cube_lut_3  = 14'b11111011110000;
        10'd825   : cube_lut_3  = 14'b11111011110010;
        10'd826   : cube_lut_3  = 14'b11111011110011;
        10'd827   : cube_lut_3  = 14'b11111011110101;
        10'd828   : cube_lut_3  = 14'b11111011110110;
        10'd829   : cube_lut_3  = 14'b11111011110111;
        10'd830   : cube_lut_3  = 14'b11111011111001;
        10'd831   : cube_lut_3  = 14'b11111011111010;
        10'd832   : cube_lut_3  = 14'b11111011111011;
        10'd833   : cube_lut_3  = 14'b11111011111101;
        10'd834   : cube_lut_3  = 14'b11111011111110;
        10'd835   : cube_lut_3  = 14'b11111100000000;
        10'd836   : cube_lut_3  = 14'b11111100000001;
        10'd837   : cube_lut_3  = 14'b11111100000010;
        10'd838   : cube_lut_3  = 14'b11111100000100;
        10'd839   : cube_lut_3  = 14'b11111100000101;
        10'd840   : cube_lut_3  = 14'b11111100000110;
        10'd841   : cube_lut_3  = 14'b11111100001000;
        10'd842   : cube_lut_3  = 14'b11111100001001;
        10'd843   : cube_lut_3  = 14'b11111100001011;
        10'd844   : cube_lut_3  = 14'b11111100001100;
        10'd845   : cube_lut_3  = 14'b11111100001101;
        10'd846   : cube_lut_3  = 14'b11111100001111;
        10'd847   : cube_lut_3  = 14'b11111100010000;
        10'd848   : cube_lut_3  = 14'b11111100010001;
        10'd849   : cube_lut_3  = 14'b11111100010011;
        10'd850   : cube_lut_3  = 14'b11111100010100;
        10'd851   : cube_lut_3  = 14'b11111100010110;
        10'd852   : cube_lut_3  = 14'b11111100010111;
        10'd853   : cube_lut_3  = 14'b11111100011000;
        10'd854   : cube_lut_3  = 14'b11111100011010;
        10'd855   : cube_lut_3  = 14'b11111100011011;
        10'd856   : cube_lut_3  = 14'b11111100011100;
        10'd857   : cube_lut_3  = 14'b11111100011110;
        10'd858   : cube_lut_3  = 14'b11111100011111;
        10'd859   : cube_lut_3  = 14'b11111100100000;
        10'd860   : cube_lut_3  = 14'b11111100100010;
        10'd861   : cube_lut_3  = 14'b11111100100011;
        10'd862   : cube_lut_3  = 14'b11111100100101;
        10'd863   : cube_lut_3  = 14'b11111100100110;
        10'd864   : cube_lut_3  = 14'b11111100100111;
        10'd865   : cube_lut_3  = 14'b11111100101001;
        10'd866   : cube_lut_3  = 14'b11111100101010;
        10'd867   : cube_lut_3  = 14'b11111100101011;
        10'd868   : cube_lut_3  = 14'b11111100101101;
        10'd869   : cube_lut_3  = 14'b11111100101110;
        10'd870   : cube_lut_3  = 14'b11111100110000;
        10'd871   : cube_lut_3  = 14'b11111100110001;
        10'd872   : cube_lut_3  = 14'b11111100110010;
        10'd873   : cube_lut_3  = 14'b11111100110100;
        10'd874   : cube_lut_3  = 14'b11111100110101;
        10'd875   : cube_lut_3  = 14'b11111100110110;
        10'd876   : cube_lut_3  = 14'b11111100111000;
        10'd877   : cube_lut_3  = 14'b11111100111001;
        10'd878   : cube_lut_3  = 14'b11111100111010;
        10'd879   : cube_lut_3  = 14'b11111100111100;
        10'd880   : cube_lut_3  = 14'b11111100111101;
        10'd881   : cube_lut_3  = 14'b11111100111111;
        10'd882   : cube_lut_3  = 14'b11111101000000;
        10'd883   : cube_lut_3  = 14'b11111101000001;
        10'd884   : cube_lut_3  = 14'b11111101000011;
        10'd885   : cube_lut_3  = 14'b11111101000100;
        10'd886   : cube_lut_3  = 14'b11111101000101;
        10'd887   : cube_lut_3  = 14'b11111101000111;
        10'd888   : cube_lut_3  = 14'b11111101001000;
        10'd889   : cube_lut_3  = 14'b11111101001001;
        10'd890   : cube_lut_3  = 14'b11111101001011;
        10'd891   : cube_lut_3  = 14'b11111101001100;
        10'd892   : cube_lut_3  = 14'b11111101001110;
        10'd893   : cube_lut_3  = 14'b11111101001111;
        10'd894   : cube_lut_3  = 14'b11111101010000;
        10'd895   : cube_lut_3  = 14'b11111101010010;
        10'd896   : cube_lut_3  = 14'b11111101010011;
        10'd897   : cube_lut_3  = 14'b11111101010100;
        10'd898   : cube_lut_3  = 14'b11111101010110;
        10'd899   : cube_lut_3  = 14'b11111101010111;
        10'd900   : cube_lut_3  = 14'b11111101011000;
        10'd901   : cube_lut_3  = 14'b11111101011010;
        10'd902   : cube_lut_3  = 14'b11111101011011;
        10'd903   : cube_lut_3  = 14'b11111101011101;
        10'd904   : cube_lut_3  = 14'b11111101011110;
        10'd905   : cube_lut_3  = 14'b11111101011111;
        10'd906   : cube_lut_3  = 14'b11111101100001;
        10'd907   : cube_lut_3  = 14'b11111101100010;
        10'd908   : cube_lut_3  = 14'b11111101100011;
        10'd909   : cube_lut_3  = 14'b11111101100101;
        10'd910   : cube_lut_3  = 14'b11111101100110;
        10'd911   : cube_lut_3  = 14'b11111101100111;
        10'd912   : cube_lut_3  = 14'b11111101101001;
        10'd913   : cube_lut_3  = 14'b11111101101010;
        10'd914   : cube_lut_3  = 14'b11111101101100;
        10'd915   : cube_lut_3  = 14'b11111101101101;
        10'd916   : cube_lut_3  = 14'b11111101101110;
        10'd917   : cube_lut_3  = 14'b11111101110000;
        10'd918   : cube_lut_3  = 14'b11111101110001;
        10'd919   : cube_lut_3  = 14'b11111101110010;
        10'd920   : cube_lut_3  = 14'b11111101110100;
        10'd921   : cube_lut_3  = 14'b11111101110101;
        10'd922   : cube_lut_3  = 14'b11111101110110;
        10'd923   : cube_lut_3  = 14'b11111101111000;
        10'd924   : cube_lut_3  = 14'b11111101111001;
        10'd925   : cube_lut_3  = 14'b11111101111010;
        10'd926   : cube_lut_3  = 14'b11111101111100;
        10'd927   : cube_lut_3  = 14'b11111101111101;
        10'd928   : cube_lut_3  = 14'b11111101111110;
        10'd929   : cube_lut_3  = 14'b11111110000000;
        10'd930   : cube_lut_3  = 14'b11111110000001;
        10'd931   : cube_lut_3  = 14'b11111110000011;
        10'd932   : cube_lut_3  = 14'b11111110000100;
        10'd933   : cube_lut_3  = 14'b11111110000101;
        10'd934   : cube_lut_3  = 14'b11111110000111;
        10'd935   : cube_lut_3  = 14'b11111110001000;
        10'd936   : cube_lut_3  = 14'b11111110001001;
        10'd937   : cube_lut_3  = 14'b11111110001011;
        10'd938   : cube_lut_3  = 14'b11111110001100;
        10'd939   : cube_lut_3  = 14'b11111110001101;
        10'd940   : cube_lut_3  = 14'b11111110001111;
        10'd941   : cube_lut_3  = 14'b11111110010000;
        10'd942   : cube_lut_3  = 14'b11111110010001;
        10'd943   : cube_lut_3  = 14'b11111110010011;
        10'd944   : cube_lut_3  = 14'b11111110010100;
        10'd945   : cube_lut_3  = 14'b11111110010101;
        10'd946   : cube_lut_3  = 14'b11111110010111;
        10'd947   : cube_lut_3  = 14'b11111110011000;
        10'd948   : cube_lut_3  = 14'b11111110011010;
        10'd949   : cube_lut_3  = 14'b11111110011011;
        10'd950   : cube_lut_3  = 14'b11111110011100;
        10'd951   : cube_lut_3  = 14'b11111110011110;
        10'd952   : cube_lut_3  = 14'b11111110011111;
        10'd953   : cube_lut_3  = 14'b11111110100000;
        10'd954   : cube_lut_3  = 14'b11111110100010;
        10'd955   : cube_lut_3  = 14'b11111110100011;
        10'd956   : cube_lut_3  = 14'b11111110100100;
        10'd957   : cube_lut_3  = 14'b11111110100110;
        10'd958   : cube_lut_3  = 14'b11111110100111;
        10'd959   : cube_lut_3  = 14'b11111110101000;
        10'd960   : cube_lut_3  = 14'b11111110101010;
        10'd961   : cube_lut_3  = 14'b11111110101011;
        10'd962   : cube_lut_3  = 14'b11111110101100;
        10'd963   : cube_lut_3  = 14'b11111110101110;
        10'd964   : cube_lut_3  = 14'b11111110101111;
        10'd965   : cube_lut_3  = 14'b11111110110000;
        10'd966   : cube_lut_3  = 14'b11111110110010;
        10'd967   : cube_lut_3  = 14'b11111110110011;
        10'd968   : cube_lut_3  = 14'b11111110110100;
        10'd969   : cube_lut_3  = 14'b11111110110110;
        10'd970   : cube_lut_3  = 14'b11111110110111;
        10'd971   : cube_lut_3  = 14'b11111110111001;
        10'd972   : cube_lut_3  = 14'b11111110111010;
        10'd973   : cube_lut_3  = 14'b11111110111011;
        10'd974   : cube_lut_3  = 14'b11111110111101;
        10'd975   : cube_lut_3  = 14'b11111110111110;
        10'd976   : cube_lut_3  = 14'b11111110111111;
        10'd977   : cube_lut_3  = 14'b11111111000001;
        10'd978   : cube_lut_3  = 14'b11111111000010;
        10'd979   : cube_lut_3  = 14'b11111111000011;
        10'd980   : cube_lut_3  = 14'b11111111000101;
        10'd981   : cube_lut_3  = 14'b11111111000110;
        10'd982   : cube_lut_3  = 14'b11111111000111;
        10'd983   : cube_lut_3  = 14'b11111111001001;
        10'd984   : cube_lut_3  = 14'b11111111001010;
        10'd985   : cube_lut_3  = 14'b11111111001011;
        10'd986   : cube_lut_3  = 14'b11111111001101;
        10'd987   : cube_lut_3  = 14'b11111111001110;
        10'd988   : cube_lut_3  = 14'b11111111001111;
        10'd989   : cube_lut_3  = 14'b11111111010001;
        10'd990   : cube_lut_3  = 14'b11111111010010;
        10'd991   : cube_lut_3  = 14'b11111111010011;
        10'd992   : cube_lut_3  = 14'b11111111010101;
        10'd993   : cube_lut_3  = 14'b11111111010110;
        10'd994   : cube_lut_3  = 14'b11111111010111;
        10'd995   : cube_lut_3  = 14'b11111111011001;
        10'd996   : cube_lut_3  = 14'b11111111011010;
        10'd997   : cube_lut_3  = 14'b11111111011011;
        10'd998   : cube_lut_3  = 14'b11111111011101;
        10'd999   : cube_lut_3  = 14'b11111111011110;
        10'd1000   : cube_lut_3 = 14'b11111111011111;
        10'd1001   : cube_lut_3 = 14'b11111111100001;
        10'd1002   : cube_lut_3 = 14'b11111111100010;
        10'd1003   : cube_lut_3 = 14'b11111111100011;
        10'd1004   : cube_lut_3 = 14'b11111111100101;
        10'd1005   : cube_lut_3 = 14'b11111111100110;
        10'd1006   : cube_lut_3 = 14'b11111111100111;
        10'd1007   : cube_lut_3 = 14'b11111111101001;
        10'd1008   : cube_lut_3 = 14'b11111111101010;
        10'd1009   : cube_lut_3 = 14'b11111111101011;
        10'd1010   : cube_lut_3 = 14'b11111111101101;
        10'd1011   : cube_lut_3 = 14'b11111111101110;
        10'd1012   : cube_lut_3 = 14'b11111111101111;
        10'd1013   : cube_lut_3 = 14'b11111111110001;
        10'd1014   : cube_lut_3 = 14'b11111111110010;
        10'd1015   : cube_lut_3 = 14'b11111111110011;
        10'd1016   : cube_lut_3 = 14'b11111111110101;
        10'd1017   : cube_lut_3 = 14'b11111111110110;
        10'd1018   : cube_lut_3 = 14'b11111111110111;
        10'd1019   : cube_lut_3 = 14'b11111111111001;
        10'd1020   : cube_lut_3 = 14'b11111111111010;
        10'd1021   : cube_lut_3 = 14'b11111111111011;
        10'd1022   : cube_lut_3 = 14'b11111111111101;
        10'd1023   : cube_lut_3 = 14'b11111111111110;
        
    endcase
end

//----------------------------------------------//
// Module Instance                              //
//----------------------------------------------//

always@(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        o_data      <= 0;
    end
    else begin
        o_data      <= o_data_nxt;
    end
end

endmodule

