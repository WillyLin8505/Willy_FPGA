// -------------------------------------------------------------------------------
// (C) Copyright. 2015
// SILICON OPTRONICS INC. ALL RIGHTS RESERVED
//
// This design is confidential and proprietary owned by Silicon Optronics Inc.
// Any distribution and modification must be authorized by a licensing agreement
// -------------------------------------------------------------------------------
// filename    : ycbcr_nominal_rng_rtl.v
// author      : Evan Tsai
//
// description : scaled & offset YCbCr(0~255) to nominal range: Y(16~235) & C(16~240) 
// -------------------------------------------------------------------------------

module ycbcr_nominal_rng(
//================================================================================
//  I/O declaratioin
//================================================================================

// output
output      [7:0]             dout_y,           //
output      [7:0]             dout_cb,          //
output      [7:0]             dout_cr,          //

// input
input       [7:0]             din_y,            //
input       [7:0]             din_cb,           //
input       [7:0]             din_cr            //
);

//================================================================================ 
//  parameter                           
//================================================================================

//================================================================================ 
//  signal declaration                             
//================================================================================
wire        [17:0]            yx879_a16;              // y*879+16
wire        [17:0]            cbx900_a16;             // cb*900+16
wire        [17:0]            crx900_a16;             // cr*900+16

//================================================================================
//  behavior description                              
//================================================================================

// YCbCr range 219
// 219/255 ~= 879(1024-128-16-1)/1024
// Yout = (Yin*879+16*1024+512)/1024
assign yx879_a16 = (din_y << 10) - (din_y << 7) - (din_y << 4) - din_y + (6'h21 << 9);
assign dout_y = (yx879_a16[17:10] > 235)? 8'd235 : yx879_a16[17:10];

// 224/255 ~= 900(1024-128+4)/1024
// Cout = (Cin*900+16*1024+512)/1024
assign cbx900_a16 = (din_cb << 10) - (din_cb << 7) + (din_cb << 2) + (6'h21 << 9);
assign dout_cb = (cbx900_a16[17:10] > 240)? 8'd240 : cbx900_a16[17:10];

assign crx900_a16 = (din_cr << 10) - (din_cr << 7) + (din_cr << 2) + (6'h21 << 9);
assign dout_cr = (crx900_a16[17:10] > 240)? 8'd240 : crx900_a16[17:10];

//================================================================================
//  module instantiation                              
//================================================================================

//================================================================================
//  function
//================================================================================
function integer log2;

input integer n;

begin
  log2 = 0;
  while(2**log2 < n) begin
    log2=log2+1;
  end
end

endfunction

//================================================================================
endmodule
